magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 990 320
<< locali >>
rect 360 25 435 55
rect 435 25 630 55
rect 435 25 465 55
rect 360 265 435 295
rect 435 265 630 295
rect 435 265 465 295
rect 360 185 435 215
rect 435 185 630 215
rect 435 185 465 215
rect 165 65 195 175
rect 180 225 255 255
rect 255 25 360 55
rect 255 25 285 255
rect 810 65 885 95
rect 810 225 885 255
rect 885 65 915 255
rect 630 105 705 135
rect 705 145 810 175
rect 705 105 735 175
rect 765 65 855 95
rect 585 185 675 215
rect 315 265 405 295
<< poly >>
rect 135 72 855 88
<< m3 >>
rect 585 0 673 320
rect 315 0 403 320
rect 585 0 673 320
rect 315 0 403 320
use JNWTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 495 160
use JNWTR_NCHDL MN1 
transform 1 0 0 0 1 80
box 0 80 495 240
use JNWTR_NCHDL MN2 
transform 1 0 0 0 1 160
box 0 160 495 320
use JNWTR_PCHDL MP0 
transform 1 0 495 0 1 0
box 495 0 990 160
use JNWTR_PCHDL MP1_DMY 
transform 1 0 495 0 1 80
box 495 80 990 240
use JNWTR_PCHDL MP2 
transform 1 0 495 0 1 160
box 495 160 990 320
use JNWTR_cut_M1M4_2x1 xcut0 
transform 1 0 585 0 1 105
box 585 105 673 139
use JNWTR_cut_M1M4_2x1 xcut1 
transform 1 0 315 0 1 105
box 315 105 403 139
use JNWTR_cut_M1M4_2x1 xcut2 
transform 1 0 315 0 1 105
box 315 105 403 139
<< labels >>
flabel locali s 765 65 855 95 0 FreeSans 400 0 0 0 C
port 1 nsew signal bidirectional
flabel locali s 585 185 675 215 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 315 265 405 295 0 FreeSans 400 0 0 0 A
port 2 nsew signal bidirectional
flabel m3 s 585 0 673 320 0 FreeSans 400 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel m3 s 315 0 403 320 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 990 320
<< end >>
