magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 648 1430
<< ppolyres >>
rect 180 -55 252 55
rect 396 -55 468 55
rect 180 55 252 165
rect 396 55 468 165
rect 180 165 252 275
rect 396 165 468 275
rect 180 275 252 385
rect 396 275 468 385
rect 180 385 252 495
rect 396 385 468 495
rect 180 495 252 605
rect 396 495 468 605
rect 180 605 252 715
rect 396 605 468 715
rect 180 715 252 825
rect 396 715 468 825
rect 180 825 252 935
rect 396 825 468 935
rect 180 935 252 1045
rect 396 935 468 1045
rect 180 1045 252 1155
rect 396 1045 468 1155
rect 180 1155 252 1265
rect 396 1155 468 1265
<< poly >>
rect -36 -55 36 55
rect 612 -55 684 55
rect -36 55 36 165
rect 612 55 684 165
rect -36 165 36 275
rect 612 165 684 275
rect -36 275 36 385
rect 612 275 684 385
rect -36 385 36 495
rect 612 385 684 495
rect -36 495 36 605
rect 612 495 684 605
rect -36 605 36 715
rect 612 605 684 715
rect -36 715 36 825
rect 612 715 684 825
rect -36 825 36 935
rect 612 825 684 935
rect -36 935 36 1045
rect 612 935 684 1045
rect -36 1045 36 1155
rect 612 1045 684 1155
rect -36 1155 36 1265
rect 612 1155 684 1265
<< xpolycontact >>
rect 180 -55 252 55
rect 396 -55 468 55
rect 180 55 252 165
rect 396 55 468 165
rect 180 1045 252 1155
rect 396 1045 468 1155
rect 180 1155 252 1265
rect 396 1155 468 1265
<< locali >>
rect 180 -55 468 55
rect 180 55 468 165
rect 180 1045 252 1155
rect 396 1045 468 1155
rect 180 1155 252 1265
rect 396 1155 468 1265
rect 180 1265 252 1375
rect 396 1265 468 1375
rect -36 1375 252 1485
rect -36 1375 252 1485
rect 396 1375 684 1485
rect 396 1375 684 1485
<< pwell >>
rect -36 -55 684 1485
<< labels >>
flabel locali s -36 1375 252 1485 0 FreeSans 400 0 0 0 N
port 1 nsew signal bidirectional
flabel locali s 396 1375 684 1485 0 FreeSans 400 0 0 0 P
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 648 1430
<< end >>
