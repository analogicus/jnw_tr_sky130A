magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 990 720
<< locali >>
rect 360 105 435 135
rect 360 265 435 295
rect 360 425 435 455
rect 360 585 435 615
rect 435 105 630 135
rect 435 265 630 295
rect 435 425 630 455
rect 435 585 630 615
rect 435 105 465 615
rect 165 65 195 655
rect 795 65 825 655
rect 135 65 225 95
rect 315 105 405 135
<< poly >>
rect 135 72 855 88
rect 135 152 855 168
rect 135 232 855 248
rect 135 312 855 328
rect 135 392 855 408
rect 135 472 855 488
rect 135 552 855 568
rect 135 632 855 648
<< m3 >>
rect 585 0 673 720
rect 315 0 403 720
rect 585 0 673 720
rect 315 0 403 720
use JNWTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 495 160
use JNWTR_NCHDL MN1 
transform 1 0 0 0 1 80
box 0 80 495 240
use JNWTR_NCHDL MN2 
transform 1 0 0 0 1 160
box 0 160 495 320
use JNWTR_NCHDL MN3 
transform 1 0 0 0 1 240
box 0 240 495 400
use JNWTR_NCHDL MN4 
transform 1 0 0 0 1 320
box 0 320 495 480
use JNWTR_NCHDL MN5 
transform 1 0 0 0 1 400
box 0 400 495 560
use JNWTR_NCHDL MN6 
transform 1 0 0 0 1 480
box 0 480 495 640
use JNWTR_NCHDL MN7 
transform 1 0 0 0 1 560
box 0 560 495 720
use JNWTR_PCHDL MP0 
transform 1 0 495 0 1 0
box 495 0 990 160
use JNWTR_PCHDL MP1 
transform 1 0 495 0 1 80
box 495 80 990 240
use JNWTR_PCHDL MP2 
transform 1 0 495 0 1 160
box 495 160 990 320
use JNWTR_PCHDL MP3 
transform 1 0 495 0 1 240
box 495 240 990 400
use JNWTR_PCHDL MP4 
transform 1 0 495 0 1 320
box 495 320 990 480
use JNWTR_PCHDL MP5 
transform 1 0 495 0 1 400
box 495 400 990 560
use JNWTR_PCHDL MP6 
transform 1 0 495 0 1 480
box 495 480 990 640
use JNWTR_PCHDL MP7 
transform 1 0 495 0 1 560
box 495 560 990 720
use JNWTR_cut_M1M4_2x1 xcut0 
transform 1 0 585 0 1 25
box 585 25 673 59
use JNWTR_cut_M1M4_2x1 xcut1 
transform 1 0 585 0 1 185
box 585 185 673 219
use JNWTR_cut_M1M4_2x1 xcut2 
transform 1 0 585 0 1 185
box 585 185 673 219
use JNWTR_cut_M1M4_2x1 xcut3 
transform 1 0 585 0 1 345
box 585 345 673 379
use JNWTR_cut_M1M4_2x1 xcut4 
transform 1 0 585 0 1 345
box 585 345 673 379
use JNWTR_cut_M1M4_2x1 xcut5 
transform 1 0 585 0 1 505
box 585 505 673 539
use JNWTR_cut_M1M4_2x1 xcut6 
transform 1 0 585 0 1 505
box 585 505 673 539
use JNWTR_cut_M1M4_2x1 xcut7 
transform 1 0 585 0 1 665
box 585 665 673 699
use JNWTR_cut_M1M4_2x1 xcut8 
transform 1 0 315 0 1 25
box 315 25 403 59
use JNWTR_cut_M1M4_2x1 xcut9 
transform 1 0 315 0 1 185
box 315 185 403 219
use JNWTR_cut_M1M4_2x1 xcut10 
transform 1 0 315 0 1 185
box 315 185 403 219
use JNWTR_cut_M1M4_2x1 xcut11 
transform 1 0 315 0 1 345
box 315 345 403 379
use JNWTR_cut_M1M4_2x1 xcut12 
transform 1 0 315 0 1 345
box 315 345 403 379
use JNWTR_cut_M1M4_2x1 xcut13 
transform 1 0 315 0 1 505
box 315 505 403 539
use JNWTR_cut_M1M4_2x1 xcut14 
transform 1 0 315 0 1 505
box 315 505 403 539
use JNWTR_cut_M1M4_2x1 xcut15 
transform 1 0 315 0 1 665
box 315 665 403 699
<< labels >>
flabel locali s 135 65 225 95 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 315 105 405 135 0 FreeSans 400 0 0 0 Y
port 2 nsew signal bidirectional
flabel m3 s 585 0 673 720 0 FreeSans 400 0 0 0 AVDD
port 3 nsew signal bidirectional
flabel m3 s 315 0 403 720 0 FreeSans 400 0 0 0 AVSS
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 990 720
<< end >>
