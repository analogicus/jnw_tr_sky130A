magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 990 400
<< locali >>
rect 180 305 255 335
rect 255 105 360 135
rect 255 105 285 335
rect 135 65 225 95
rect 135 145 225 175
rect 315 345 405 375
<< m3 >>
rect 585 0 673 400
rect 315 0 403 400
rect 585 0 673 400
rect 315 0 403 400
use JNWTR_NRX1_CV XA1 
transform 1 0 0 0 1 0
box 0 0 990 240
use JNWTR_IVX1_CV XA2 
transform 1 0 0 0 1 240
box 0 240 990 400
<< labels >>
flabel locali s 135 65 225 95 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 135 145 225 175 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel locali s 315 345 405 375 0 FreeSans 400 0 0 0 Y
port 3 nsew signal bidirectional
flabel m3 s 585 0 673 400 0 FreeSans 400 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel m3 s 315 0 403 400 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 990 400
<< end >>
