magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 88 34
<< m3 >>
rect 0 0 88 34
<< v3 >>
rect 6 3 34 31
rect 54 3 82 31
<< m4 >>
rect 0 0 88 34
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 88 34
<< end >>
