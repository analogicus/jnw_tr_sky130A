magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 2632 2118
<< locali >>
rect 8 8 2624 64
rect 64 8 2568 64
rect 8 8 2624 64
rect 64 2054 2568 2110
rect 8 2054 2624 2110
rect 8 64 64 2054
rect 8 8 64 2110
rect 2568 64 2624 2054
rect 2568 8 2624 2110
rect 8 8 2624 64
rect 2036 1719 2324 1829
rect 308 1719 596 1829
<< ptapc >>
rect 76 16 116 56
rect 116 16 156 56
rect 156 16 196 56
rect 196 16 236 56
rect 236 16 276 56
rect 276 16 316 56
rect 316 16 356 56
rect 356 16 396 56
rect 396 16 436 56
rect 436 16 476 56
rect 476 16 516 56
rect 516 16 556 56
rect 556 16 596 56
rect 596 16 636 56
rect 636 16 676 56
rect 676 16 716 56
rect 716 16 756 56
rect 756 16 796 56
rect 796 16 836 56
rect 836 16 876 56
rect 876 16 916 56
rect 916 16 956 56
rect 956 16 996 56
rect 996 16 1036 56
rect 1036 16 1076 56
rect 1076 16 1116 56
rect 1116 16 1156 56
rect 1156 16 1196 56
rect 1196 16 1236 56
rect 1236 16 1276 56
rect 1276 16 1316 56
rect 1316 16 1356 56
rect 1356 16 1396 56
rect 1396 16 1436 56
rect 1436 16 1476 56
rect 1476 16 1516 56
rect 1516 16 1556 56
rect 1556 16 1596 56
rect 1596 16 1636 56
rect 1636 16 1676 56
rect 1676 16 1716 56
rect 1716 16 1756 56
rect 1756 16 1796 56
rect 1796 16 1836 56
rect 1836 16 1876 56
rect 1876 16 1916 56
rect 1916 16 1956 56
rect 1956 16 1996 56
rect 1996 16 2036 56
rect 2036 16 2076 56
rect 2076 16 2116 56
rect 2116 16 2156 56
rect 2156 16 2196 56
rect 2196 16 2236 56
rect 2236 16 2276 56
rect 2276 16 2316 56
rect 2316 16 2356 56
rect 2356 16 2396 56
rect 2396 16 2436 56
rect 2436 16 2476 56
rect 2476 16 2516 56
rect 2516 16 2556 56
rect 76 2062 116 2102
rect 116 2062 156 2102
rect 156 2062 196 2102
rect 196 2062 236 2102
rect 236 2062 276 2102
rect 276 2062 316 2102
rect 316 2062 356 2102
rect 356 2062 396 2102
rect 396 2062 436 2102
rect 436 2062 476 2102
rect 476 2062 516 2102
rect 516 2062 556 2102
rect 556 2062 596 2102
rect 596 2062 636 2102
rect 636 2062 676 2102
rect 676 2062 716 2102
rect 716 2062 756 2102
rect 756 2062 796 2102
rect 796 2062 836 2102
rect 836 2062 876 2102
rect 876 2062 916 2102
rect 916 2062 956 2102
rect 956 2062 996 2102
rect 996 2062 1036 2102
rect 1036 2062 1076 2102
rect 1076 2062 1116 2102
rect 1116 2062 1156 2102
rect 1156 2062 1196 2102
rect 1196 2062 1236 2102
rect 1236 2062 1276 2102
rect 1276 2062 1316 2102
rect 1316 2062 1356 2102
rect 1356 2062 1396 2102
rect 1396 2062 1436 2102
rect 1436 2062 1476 2102
rect 1476 2062 1516 2102
rect 1516 2062 1556 2102
rect 1556 2062 1596 2102
rect 1596 2062 1636 2102
rect 1636 2062 1676 2102
rect 1676 2062 1716 2102
rect 1716 2062 1756 2102
rect 1756 2062 1796 2102
rect 1796 2062 1836 2102
rect 1836 2062 1876 2102
rect 1876 2062 1916 2102
rect 1916 2062 1956 2102
rect 1956 2062 1996 2102
rect 1996 2062 2036 2102
rect 2036 2062 2076 2102
rect 2076 2062 2116 2102
rect 2116 2062 2156 2102
rect 2156 2062 2196 2102
rect 2196 2062 2236 2102
rect 2236 2062 2276 2102
rect 2276 2062 2316 2102
rect 2316 2062 2356 2102
rect 2356 2062 2396 2102
rect 2396 2062 2436 2102
rect 2436 2062 2476 2102
rect 2476 2062 2516 2102
rect 2516 2062 2556 2102
rect 16 79 56 119
rect 16 119 56 159
rect 16 159 56 199
rect 16 199 56 239
rect 16 239 56 279
rect 16 279 56 319
rect 16 319 56 359
rect 16 359 56 399
rect 16 399 56 439
rect 16 439 56 479
rect 16 479 56 519
rect 16 519 56 559
rect 16 559 56 599
rect 16 599 56 639
rect 16 639 56 679
rect 16 679 56 719
rect 16 719 56 759
rect 16 759 56 799
rect 16 799 56 839
rect 16 839 56 879
rect 16 879 56 919
rect 16 919 56 959
rect 16 959 56 999
rect 16 999 56 1039
rect 16 1039 56 1079
rect 16 1079 56 1119
rect 16 1119 56 1159
rect 16 1159 56 1199
rect 16 1199 56 1239
rect 16 1239 56 1279
rect 16 1279 56 1319
rect 16 1319 56 1359
rect 16 1359 56 1399
rect 16 1399 56 1439
rect 16 1439 56 1479
rect 16 1479 56 1519
rect 16 1519 56 1559
rect 16 1559 56 1599
rect 16 1599 56 1639
rect 16 1639 56 1679
rect 16 1679 56 1719
rect 16 1719 56 1759
rect 16 1759 56 1799
rect 16 1799 56 1839
rect 16 1839 56 1879
rect 16 1879 56 1919
rect 16 1919 56 1959
rect 16 1959 56 1999
rect 16 1999 56 2039
rect 2576 79 2616 119
rect 2576 119 2616 159
rect 2576 159 2616 199
rect 2576 199 2616 239
rect 2576 239 2616 279
rect 2576 279 2616 319
rect 2576 319 2616 359
rect 2576 359 2616 399
rect 2576 399 2616 439
rect 2576 439 2616 479
rect 2576 479 2616 519
rect 2576 519 2616 559
rect 2576 559 2616 599
rect 2576 599 2616 639
rect 2576 639 2616 679
rect 2576 679 2616 719
rect 2576 719 2616 759
rect 2576 759 2616 799
rect 2576 799 2616 839
rect 2576 839 2616 879
rect 2576 879 2616 919
rect 2576 919 2616 959
rect 2576 959 2616 999
rect 2576 999 2616 1039
rect 2576 1039 2616 1079
rect 2576 1079 2616 1119
rect 2576 1119 2616 1159
rect 2576 1159 2616 1199
rect 2576 1199 2616 1239
rect 2576 1239 2616 1279
rect 2576 1279 2616 1319
rect 2576 1319 2616 1359
rect 2576 1359 2616 1399
rect 2576 1399 2616 1439
rect 2576 1439 2616 1479
rect 2576 1479 2616 1519
rect 2576 1519 2616 1559
rect 2576 1559 2616 1599
rect 2576 1599 2616 1639
rect 2576 1639 2616 1679
rect 2576 1679 2616 1719
rect 2576 1719 2616 1759
rect 2576 1759 2616 1799
rect 2576 1799 2616 1839
rect 2576 1839 2616 1879
rect 2576 1879 2616 1919
rect 2576 1919 2616 1959
rect 2576 1959 2616 1999
rect 2576 1999 2616 2039
<< ptap >>
rect 0 0 2632 72
rect 0 2046 2632 2118
rect 0 0 72 2118
rect 2560 0 2632 2118
use JNWTR_RES8 XA1 
transform 1 0 344 0 1 344
box 344 344 2288 1774
<< labels >>
flabel locali s 8 8 2624 64 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 2036 1719 2324 1829 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel locali s 308 1719 596 1829 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2632 2118
<< end >>
