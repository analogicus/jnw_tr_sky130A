magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1260 264
<< locali >>
rect 216 161 300 191
rect 300 29 432 59
rect 300 29 330 191
rect 432 29 516 59
rect 516 29 828 59
rect 516 29 546 59
rect 432 205 516 235
rect 516 205 828 235
rect 516 205 546 235
rect 162 73 270 103
rect 378 205 486 235
<< poly >>
rect 162 79 1098 97
rect 162 167 1098 185
<< m3 >>
rect 774 0 874 264
rect 378 0 478 264
rect 774 0 874 264
rect 378 0 478 264
use JNWTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 630 176
use JNWTR_NCHDL MN1 
transform 1 0 0 0 1 88
box 0 88 630 264
use JNWTR_PCHDL MP0 
transform 1 0 630 0 1 0
box 630 0 1260 176
use JNWTR_PCHDL MP1 
transform 1 0 630 0 1 88
box 630 88 1260 264
use JNWTR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 117
box 774 117 874 155
use JNWTR_cut_M1M4_2x1 xcut1 
transform 1 0 774 0 1 117
box 774 117 874 155
use JNWTR_cut_M1M4_2x1 xcut2 
transform 1 0 378 0 1 117
box 378 117 478 155
use JNWTR_cut_M1M4_2x1 xcut3 
transform 1 0 378 0 1 117
box 378 117 478 155
<< labels >>
flabel locali s 162 73 270 103 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 378 205 486 235 0 FreeSans 400 0 0 0 Y
port 2 nsew signal bidirectional
flabel m3 s 774 0 874 264 0 FreeSans 400 0 0 0 AVDD
port 3 nsew signal bidirectional
flabel m3 s 378 0 478 264 0 FreeSans 400 0 0 0 AVSS
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 264
<< end >>
