magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 990 480
<< locali >>
rect 345 265 375 375
rect 615 105 645 215
rect 360 185 435 215
rect 435 425 630 455
rect 435 185 465 455
rect 75 385 180 415
rect 75 135 345 165
rect 75 135 105 415
rect 315 105 360 135
rect 360 105 495 135
rect 495 265 630 295
rect 495 105 525 295
rect 135 65 225 95
rect 135 225 225 255
rect 315 185 405 215
<< poly >>
rect 135 72 855 88
rect 135 232 855 248
rect 135 392 855 408
<< m3 >>
rect 585 0 673 480
rect 315 0 403 480
rect 585 0 673 480
rect 315 0 403 480
use JNWTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 495 160
use JNWTR_NCHDL MN2 
transform 1 0 0 0 1 160
box 0 160 495 320
use JNWTR_NCHDL MN1 
transform 1 0 0 0 1 320
box 0 320 495 480
use JNWTR_PCHDL MP1 
transform 1 0 495 0 1 0
box 495 0 990 160
use JNWTR_PCHDL MP0 
transform 1 0 495 0 1 160
box 495 160 990 320
use JNWTR_PCHDL MP2 
transform 1 0 495 0 1 320
box 495 320 990 480
use JNWTR_cut_M1M4_2x1 xcut0 
transform 1 0 585 0 1 25
box 585 25 673 59
use JNWTR_cut_M1M4_2x1 xcut1 
transform 1 0 585 0 1 345
box 585 345 673 379
use JNWTR_cut_M1M4_2x1 xcut2 
transform 1 0 315 0 1 25
box 315 25 403 59
use JNWTR_cut_M1M4_2x1 xcut3 
transform 1 0 315 0 1 425
box 315 425 403 459
<< labels >>
flabel locali s 135 65 225 95 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 135 225 225 255 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 315 185 405 215 0 FreeSans 400 0 0 0 Q
port 3 nsew signal bidirectional
flabel m3 s 585 0 673 480 0 FreeSans 400 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel m3 s 315 0 403 480 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 990 480
<< end >>
