magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 60 0 1200 1140
<< m3 >>
rect 500 0 930 40
rect 330 600 500 640
rect 330 0 500 40
rect 500 600 930 640
rect 500 0 540 640
rect 60 0 600 50
<< m4 >>
rect 500 0 930 40
rect 330 600 500 640
rect 330 0 500 40
rect 500 600 930 640
rect 500 0 540 640
rect 60 0 600 50
use JNWTR_CAPX1 XA1 
transform 1 0 60 0 1 0
box 60 0 600 540
use JNWTR_CAPX1 XA2 
transform 1 0 60 0 1 600
box 60 600 600 1140
use JNWTR_CAPX1 XB1 
transform 1 0 660 0 1 0
box 660 0 1200 540
use JNWTR_CAPX1 XB2 
transform 1 0 660 0 1 600
box 660 600 1200 1140
<< labels >>
flabel m3 s 60 0 600 50 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel m4 s 60 0 600 50 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 60 0 1200 1140
<< end >>
