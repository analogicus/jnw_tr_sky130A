magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 720 176
<< ndiff >>
rect 378 22 486 66
rect 378 66 486 110
rect 378 110 486 154
<< ptap >>
rect -54 -22 54 22
rect -54 22 54 66
rect -54 66 54 110
rect -54 110 54 154
rect -54 154 54 198
<< poly >>
rect 162 -9 522 9
rect 162 79 522 97
rect 162 167 522 185
rect 162 66 270 110
<< locali >>
rect 162 73 270 103
rect -54 -22 54 22
rect -54 22 54 66
rect 378 29 486 59
rect 378 29 486 59
rect -54 66 54 110
rect -54 66 54 110
rect 162 73 270 103
rect -54 110 54 154
rect 378 117 486 147
rect 378 117 486 147
rect -54 154 54 198
<< pcontact >>
rect 174 77 198 88
rect 174 88 198 99
rect 198 77 234 88
rect 198 88 234 99
rect 234 77 258 88
rect 234 88 258 99
<< ptapc >>
rect -18 22 18 66
rect -18 110 18 154
<< ndcontact >>
rect 390 33 414 44
rect 390 44 414 55
rect 414 33 450 44
rect 414 44 450 55
rect 450 33 474 44
rect 450 44 474 55
rect 390 121 414 132
rect 390 132 414 143
rect 414 121 450 132
rect 414 132 450 143
rect 450 121 474 132
rect 450 132 474 143
<< pwell >>
rect -90 -66 630 242
<< labels >>
flabel locali s 162 73 270 103 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 378 29 486 59 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s -54 66 54 110 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 378 117 486 147 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 720 176
<< end >>
