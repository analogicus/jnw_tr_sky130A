magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1768 2118
<< locali >>
rect 8 8 1760 64
rect 64 8 1704 64
rect 8 8 1760 64
rect 64 2054 1704 2110
rect 8 2054 1760 2110
rect 8 64 64 2054
rect 8 8 64 2110
rect 1704 64 1760 2054
rect 1704 8 1760 2110
rect 8 8 1760 64
rect 1172 1719 1460 1829
rect 308 1719 596 1829
<< ptapc >>
rect 84 16 124 56
rect 124 16 164 56
rect 164 16 204 56
rect 204 16 244 56
rect 244 16 284 56
rect 284 16 324 56
rect 324 16 364 56
rect 364 16 404 56
rect 404 16 444 56
rect 444 16 484 56
rect 484 16 524 56
rect 524 16 564 56
rect 564 16 604 56
rect 604 16 644 56
rect 644 16 684 56
rect 684 16 724 56
rect 724 16 764 56
rect 764 16 804 56
rect 804 16 844 56
rect 844 16 884 56
rect 884 16 924 56
rect 924 16 964 56
rect 964 16 1004 56
rect 1004 16 1044 56
rect 1044 16 1084 56
rect 1084 16 1124 56
rect 1124 16 1164 56
rect 1164 16 1204 56
rect 1204 16 1244 56
rect 1244 16 1284 56
rect 1284 16 1324 56
rect 1324 16 1364 56
rect 1364 16 1404 56
rect 1404 16 1444 56
rect 1444 16 1484 56
rect 1484 16 1524 56
rect 1524 16 1564 56
rect 1564 16 1604 56
rect 1604 16 1644 56
rect 1644 16 1684 56
rect 84 2062 124 2102
rect 124 2062 164 2102
rect 164 2062 204 2102
rect 204 2062 244 2102
rect 244 2062 284 2102
rect 284 2062 324 2102
rect 324 2062 364 2102
rect 364 2062 404 2102
rect 404 2062 444 2102
rect 444 2062 484 2102
rect 484 2062 524 2102
rect 524 2062 564 2102
rect 564 2062 604 2102
rect 604 2062 644 2102
rect 644 2062 684 2102
rect 684 2062 724 2102
rect 724 2062 764 2102
rect 764 2062 804 2102
rect 804 2062 844 2102
rect 844 2062 884 2102
rect 884 2062 924 2102
rect 924 2062 964 2102
rect 964 2062 1004 2102
rect 1004 2062 1044 2102
rect 1044 2062 1084 2102
rect 1084 2062 1124 2102
rect 1124 2062 1164 2102
rect 1164 2062 1204 2102
rect 1204 2062 1244 2102
rect 1244 2062 1284 2102
rect 1284 2062 1324 2102
rect 1324 2062 1364 2102
rect 1364 2062 1404 2102
rect 1404 2062 1444 2102
rect 1444 2062 1484 2102
rect 1484 2062 1524 2102
rect 1524 2062 1564 2102
rect 1564 2062 1604 2102
rect 1604 2062 1644 2102
rect 1644 2062 1684 2102
rect 16 79 56 119
rect 16 119 56 159
rect 16 159 56 199
rect 16 199 56 239
rect 16 239 56 279
rect 16 279 56 319
rect 16 319 56 359
rect 16 359 56 399
rect 16 399 56 439
rect 16 439 56 479
rect 16 479 56 519
rect 16 519 56 559
rect 16 559 56 599
rect 16 599 56 639
rect 16 639 56 679
rect 16 679 56 719
rect 16 719 56 759
rect 16 759 56 799
rect 16 799 56 839
rect 16 839 56 879
rect 16 879 56 919
rect 16 919 56 959
rect 16 959 56 999
rect 16 999 56 1039
rect 16 1039 56 1079
rect 16 1079 56 1119
rect 16 1119 56 1159
rect 16 1159 56 1199
rect 16 1199 56 1239
rect 16 1239 56 1279
rect 16 1279 56 1319
rect 16 1319 56 1359
rect 16 1359 56 1399
rect 16 1399 56 1439
rect 16 1439 56 1479
rect 16 1479 56 1519
rect 16 1519 56 1559
rect 16 1559 56 1599
rect 16 1599 56 1639
rect 16 1639 56 1679
rect 16 1679 56 1719
rect 16 1719 56 1759
rect 16 1759 56 1799
rect 16 1799 56 1839
rect 16 1839 56 1879
rect 16 1879 56 1919
rect 16 1919 56 1959
rect 16 1959 56 1999
rect 16 1999 56 2039
rect 1712 79 1752 119
rect 1712 119 1752 159
rect 1712 159 1752 199
rect 1712 199 1752 239
rect 1712 239 1752 279
rect 1712 279 1752 319
rect 1712 319 1752 359
rect 1712 359 1752 399
rect 1712 399 1752 439
rect 1712 439 1752 479
rect 1712 479 1752 519
rect 1712 519 1752 559
rect 1712 559 1752 599
rect 1712 599 1752 639
rect 1712 639 1752 679
rect 1712 679 1752 719
rect 1712 719 1752 759
rect 1712 759 1752 799
rect 1712 799 1752 839
rect 1712 839 1752 879
rect 1712 879 1752 919
rect 1712 919 1752 959
rect 1712 959 1752 999
rect 1712 999 1752 1039
rect 1712 1039 1752 1079
rect 1712 1079 1752 1119
rect 1712 1119 1752 1159
rect 1712 1159 1752 1199
rect 1712 1199 1752 1239
rect 1712 1239 1752 1279
rect 1712 1279 1752 1319
rect 1712 1319 1752 1359
rect 1712 1359 1752 1399
rect 1712 1399 1752 1439
rect 1712 1439 1752 1479
rect 1712 1479 1752 1519
rect 1712 1519 1752 1559
rect 1712 1559 1752 1599
rect 1712 1599 1752 1639
rect 1712 1639 1752 1679
rect 1712 1679 1752 1719
rect 1712 1719 1752 1759
rect 1712 1759 1752 1799
rect 1712 1799 1752 1839
rect 1712 1839 1752 1879
rect 1712 1879 1752 1919
rect 1712 1919 1752 1959
rect 1712 1959 1752 1999
rect 1712 1999 1752 2039
<< ptap >>
rect 0 0 1768 72
rect 0 2046 1768 2118
rect 0 0 72 2118
rect 1696 0 1768 2118
use JNWTR_RES4 XA1 
transform 1 0 344 0 1 344
box 344 344 1424 1774
<< labels >>
flabel locali s 8 8 1760 64 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 1172 1719 1460 1829 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel locali s 308 1719 596 1829 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1768 2118
<< end >>
