magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1260 264
<< locali >>
rect 432 205 516 235
rect 516 117 828 147
rect 516 117 546 235
rect 417 117 447 147
rect 162 73 270 103
rect 162 161 270 191
rect 378 205 486 235
<< poly >>
rect 162 79 1098 97
rect 162 167 1098 185
<< m3 >>
rect 774 0 874 264
rect 378 0 478 264
rect 774 0 874 264
rect 378 0 478 264
use JNWTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 630 176
use JNWTR_NCHDL MN1 
transform 1 0 0 0 1 88
box 0 88 630 264
use JNWTR_PCHDL MP0 
transform 1 0 630 0 1 0
box 630 0 1260 176
use JNWTR_PCHDL MP1 
transform 1 0 630 0 1 88
box 630 88 1260 264
use JNWTR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 29
box 774 29 874 67
use JNWTR_cut_M1M4_2x1 xcut1 
transform 1 0 774 0 1 205
box 774 205 874 243
use JNWTR_cut_M1M4_2x1 xcut2 
transform 1 0 378 0 1 29
box 378 29 478 67
<< labels >>
flabel locali s 162 73 270 103 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 162 161 270 191 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel locali s 378 205 486 235 0 FreeSans 400 0 0 0 Y
port 3 nsew signal bidirectional
flabel m3 s 774 0 874 264 0 FreeSans 400 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel m3 s 378 0 478 264 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 264
<< end >>
