magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 940 1720
<< locali >>
rect 8 8 932 64
rect 64 8 876 64
rect 8 8 932 64
rect 64 1656 876 1712
rect 8 1656 932 1712
rect 8 64 64 1656
rect 8 8 64 1712
rect 876 64 932 1656
rect 876 8 932 1712
rect 8 8 932 64
rect 614 1460 758 1580
rect 182 1460 326 1580
<< ptapc >>
rect 90 16 130 56
rect 130 16 170 56
rect 170 16 210 56
rect 210 16 250 56
rect 250 16 290 56
rect 290 16 330 56
rect 330 16 370 56
rect 370 16 410 56
rect 410 16 450 56
rect 450 16 490 56
rect 490 16 530 56
rect 530 16 570 56
rect 570 16 610 56
rect 610 16 650 56
rect 650 16 690 56
rect 690 16 730 56
rect 730 16 770 56
rect 770 16 810 56
rect 810 16 850 56
rect 90 1664 130 1704
rect 130 1664 170 1704
rect 170 1664 210 1704
rect 210 1664 250 1704
rect 250 1664 290 1704
rect 290 1664 330 1704
rect 330 1664 370 1704
rect 370 1664 410 1704
rect 410 1664 450 1704
rect 450 1664 490 1704
rect 490 1664 530 1704
rect 530 1664 570 1704
rect 570 1664 610 1704
rect 610 1664 650 1704
rect 650 1664 690 1704
rect 690 1664 730 1704
rect 730 1664 770 1704
rect 770 1664 810 1704
rect 810 1664 850 1704
rect 16 80 56 120
rect 16 120 56 160
rect 16 160 56 200
rect 16 200 56 240
rect 16 240 56 280
rect 16 280 56 320
rect 16 320 56 360
rect 16 360 56 400
rect 16 400 56 440
rect 16 440 56 480
rect 16 480 56 520
rect 16 520 56 560
rect 16 560 56 600
rect 16 600 56 640
rect 16 640 56 680
rect 16 680 56 720
rect 16 720 56 760
rect 16 760 56 800
rect 16 800 56 840
rect 16 840 56 880
rect 16 880 56 920
rect 16 920 56 960
rect 16 960 56 1000
rect 16 1000 56 1040
rect 16 1040 56 1080
rect 16 1080 56 1120
rect 16 1120 56 1160
rect 16 1160 56 1200
rect 16 1200 56 1240
rect 16 1240 56 1280
rect 16 1280 56 1320
rect 16 1320 56 1360
rect 16 1360 56 1400
rect 16 1400 56 1440
rect 16 1440 56 1480
rect 16 1480 56 1520
rect 16 1520 56 1560
rect 16 1560 56 1600
rect 16 1600 56 1640
rect 884 80 924 120
rect 884 120 924 160
rect 884 160 924 200
rect 884 200 924 240
rect 884 240 924 280
rect 884 280 924 320
rect 884 320 924 360
rect 884 360 924 400
rect 884 400 924 440
rect 884 440 924 480
rect 884 480 924 520
rect 884 520 924 560
rect 884 560 924 600
rect 884 600 924 640
rect 884 640 924 680
rect 884 680 924 720
rect 884 720 924 760
rect 884 760 924 800
rect 884 800 924 840
rect 884 840 924 880
rect 884 880 924 920
rect 884 920 924 960
rect 884 960 924 1000
rect 884 1000 924 1040
rect 884 1040 924 1080
rect 884 1080 924 1120
rect 884 1120 924 1160
rect 884 1160 924 1200
rect 884 1200 924 1240
rect 884 1240 924 1280
rect 884 1280 924 1320
rect 884 1320 924 1360
rect 884 1360 924 1400
rect 884 1400 924 1440
rect 884 1440 924 1480
rect 884 1480 924 1520
rect 884 1520 924 1560
rect 884 1560 924 1600
rect 884 1600 924 1640
<< ptap >>
rect 0 0 940 72
rect 0 1648 940 1720
rect 0 0 72 1720
rect 868 0 940 1720
use JNWTR_RES4 XA1 
transform 1 0 200 0 1 200
box 200 200 740 1520
<< labels >>
flabel locali s 8 8 932 64 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 614 1460 758 1580 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel locali s 182 1460 326 1580 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 940 1720
<< end >>
