

.subckt TGX2_CV A C B AVDD AVSS
MN0 AVSS C CN AVSS NCHDL
MN1 B C A AVSS NCHDL
MN1b B C A AVSS NCHDL

MP0 AVDD C CN AVDD PCHDL
MP1 B CN A AVDD PCHDL
MP1b B CN A AVDD PCHDL

.ends

.subckt DFTRIX1_CV D CK C CN Y AVDD AVSS
XA3 AVDD AVSS TAPCELLB_CV
XA2 D CK C NC QN AVDD AVSS DFRNQNX1_CV
XA0 QN C CN Y AVDD AVSS IVTRIX1_CV
.ends


.SUBCKT CKDIV2 AVDD AVSS CKI CKO CKO50DC RN
XA12v AVDD AVSS TAPCELLB_CV
XA1 CKI CKIB AVDD AVSS BFX1_CV
XA2 CKIB CKIN AVDD AVSS  IVX1_CV
XA4  QNI CKIN RN CKO50DC QN AVDD AVSS DFRNQNX1_CV
XA3 CKO50DC QNI AVDD AVSS  IVX1_CV
XA5 CKO50DC CKI CKO AVDD AVSS ANX1_CV

.ENDS

.subckt RG12TRIX1_CV D<11> D<10> D<9> D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0> CK C CN
+ Y<11> Y<10> Y<9> Y<8> Y<7> Y<6> Y<5> Y<4> Y<3> Y<2> Y<1> Y<0> AVDD AVSS
XA0 D<11> CK C CN Y<11> AVDD AVSS DFTRIX1_CV
XB1 D<10> CK C CN Y<10> AVDD AVSS DFTRIX1_CV
XC2 D<9> CK C CN Y<9> AVDD AVSS DFTRIX1_CV
XD3 D<8> CK C CN Y<8> AVDD AVSS DFTRIX1_CV
XE4 D<7> CK C CN Y<7> AVDD AVSS DFTRIX1_CV
XF5 D<6> CK C CN Y<6> AVDD AVSS DFTRIX1_CV
XG6 D<5> CK C CN Y<5> AVDD AVSS DFTRIX1_CV
XH7 D<4> CK C CN Y<4> AVDD AVSS DFTRIX1_CV
XI8 D<3> CK C CN Y<3> AVDD AVSS DFTRIX1_CV
XJ9 D<2> CK C CN Y<2> AVDD AVSS DFTRIX1_CV
XK10 D<1> CK C CN Y<1> AVDD AVSS DFTRIX1_CV
XL11 D<0> CK C CN Y<0> AVDD AVSS DFTRIX1_CV
.ends


.subckt TOP AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA1 Y1 AVDD AVSS TIEH_CV
XA2 Y2 AVDD AVSS TIEL_CV
XB0 AVDD AVSS TAPCELLB_CV
XB3 A3 Y3 AVDD AVSS IVX1_CV
XB4 A4 Y4 AVDD AVSS IVX2_CV
XB5 A5 Y5 AVDD AVSS IVX4_CV
XB6 A6 Y6 AVDD AVSS IVX8_CV
XC0 AVDD AVSS TAPCELLB_CV
XC7 A7 Y7 AVDD AVSS BFX1_CV
XD0 AVDD AVSS TAPCELLB_CV
XD8 A8 B8 Y8 AVDD AVSS NRX1_CV
XD9 A9 B9 Y9 AVDD AVSS NDX1_CV
XD10 A10 B10 Y10 AVDD AVSS ORX1_CV
XD11 A11 B11 Y11 AVDD AVSS ANX1_CV
XE0 AVDD AVSS TAPCELLB_CV
XE12 A12 Y12 AVDD AVSS SCX1_CV
XF0 AVDD AVSS TAPCELLB_CV
XF13 A13 Y13 V13 AVDD AVSS SWX2_CV
XF14 A14 Y14 V14 AVDD AVSS SWX4_CV
XF15 A15 Y15 V15 AVDD AVSS TGPD_CV
XG0 AVDD AVSS TAPCELLB_CV
XG1 A16 C16 B16 AVDD AVSS TGX2_CV
XH1 P17 N17 AVSS RPPO2 xoffset=4
XI1 P18 N18 AVSS RPPO4 xoffset=4
XJ1 P19 N19 AVSS RPPO8 xoffset=4
XK1 P20 N20 AVSS RPPO16 xoffset=4
.ends
