magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1260 2112
<< locali >>
rect 828 293 912 323
rect 912 483 1020 513
rect 912 293 942 513
rect 990 513 1044 543
rect 828 557 912 587
rect 912 777 1044 807
rect 912 1833 1044 1863
rect 912 557 942 1863
rect 216 1041 300 1071
rect 300 557 432 587
rect 300 557 330 1071
rect 240 1451 300 1481
rect 300 557 432 587
rect 300 557 330 1481
rect 216 1481 270 1511
rect 432 821 516 851
rect 432 1085 516 1115
rect 516 821 546 1115
rect 216 2009 300 2039
rect 300 1877 432 1907
rect 300 1877 330 2039
rect 990 689 1098 719
rect 162 249 270 279
rect 378 2053 486 2083
rect 378 1877 486 1907
rect 162 1657 270 1687
<< m1 >>
rect 1044 1041 1128 1071
rect 1044 1481 1128 1511
rect 828 293 1128 323
rect 1128 293 1158 1511
rect 240 747 300 777
rect 300 381 432 411
rect 300 381 330 777
rect 216 777 270 807
rect 432 1525 516 1555
rect 432 1877 516 1907
rect 516 1525 546 1907
rect 216 1217 300 1247
rect 300 1085 432 1115
rect 300 1085 330 1247
rect 828 1261 912 1291
rect 912 953 1044 983
rect 912 1393 1044 1423
rect 912 953 942 1423
rect 828 2053 912 2083
rect 912 1745 1044 1775
rect 912 1745 942 2083
rect 102 337 216 367
rect 102 1657 216 1687
rect 102 337 132 1687
<< m2 >>
rect 216 1833 302 1871
rect 302 1481 1044 1519
rect 302 1481 340 1871
<< m3 >>
rect 774 0 874 2112
rect 378 0 478 2112
rect 774 0 874 2112
rect 378 0 478 2112
use JNWTR_TAPCELLB_CV XA0 
transform 1 0 0 0 1 0
box 0 0 1260 176
use JNWTR_NDX1_CV XA1 
transform 1 0 0 0 1 176
box 0 176 1260 440
use JNWTR_IVX1_CV XA2 
transform 1 0 0 0 1 440
box 0 440 1260 616
use JNWTR_IVTRIX1_CV XA3 
transform 1 0 0 0 1 616
box 0 616 1260 880
use JNWTR_IVTRIX1_CV XA4 
transform 1 0 0 0 1 880
box 0 880 1260 1144
use JNWTR_IVX1_CV XA5 
transform 1 0 0 0 1 1144
box 0 1144 1260 1320
use JNWTR_IVTRIX1_CV XA6 
transform 1 0 0 0 1 1320
box 0 1320 1260 1584
use JNWTR_NDTRIX1_CV XA7 
transform 1 0 0 0 1 1584
box 0 1584 1260 1936
use JNWTR_IVX1_CV XA8 
transform 1 0 0 0 1 1936
box 0 1936 1260 2112
use JNWTR_cut_M1M2_2x1 xcut0 
transform 1 0 990 0 1 1041
box 990 1041 1082 1075
use JNWTR_cut_M1M2_2x1 xcut1 
transform 1 0 990 0 1 1481
box 990 1481 1082 1515
use JNWTR_cut_M1M2_2x1 xcut2 
transform 1 0 774 0 1 293
box 774 293 866 327
use JNWTR_cut_M1M2_2x1 xcut3 
transform 1 0 162 0 1 777
box 162 777 254 811
use JNWTR_cut_M1M2_2x1 xcut4 
transform 1 0 378 0 1 381
box 378 381 470 415
use JNWTR_cut_M1M3_2x1 xcut5 
transform 1 0 162 0 1 1833
box 162 1833 262 1871
use JNWTR_cut_M1M3_2x1 xcut6 
transform 1 0 990 0 1 1481
box 990 1481 1090 1519
use JNWTR_cut_M1M2_2x1 xcut7 
transform 1 0 378 0 1 1525
box 378 1525 470 1559
use JNWTR_cut_M1M2_2x1 xcut8 
transform 1 0 378 0 1 1877
box 378 1877 470 1911
use JNWTR_cut_M1M2_2x1 xcut9 
transform 1 0 162 0 1 1217
box 162 1217 254 1251
use JNWTR_cut_M1M2_2x1 xcut10 
transform 1 0 378 0 1 1085
box 378 1085 470 1119
use JNWTR_cut_M1M2_2x1 xcut11 
transform 1 0 774 0 1 1261
box 774 1261 866 1295
use JNWTR_cut_M1M2_2x1 xcut12 
transform 1 0 990 0 1 953
box 990 953 1082 987
use JNWTR_cut_M1M2_2x1 xcut13 
transform 1 0 990 0 1 1393
box 990 1393 1082 1427
use JNWTR_cut_M1M2_2x1 xcut14 
transform 1 0 774 0 1 2053
box 774 2053 866 2087
use JNWTR_cut_M1M2_2x1 xcut15 
transform 1 0 990 0 1 1745
box 990 1745 1082 1779
use JNWTR_cut_M1M2_2x1 xcut16 
transform 1 0 162 0 1 337
box 162 337 254 371
use JNWTR_cut_M1M2_2x1 xcut17 
transform 1 0 162 0 1 1657
box 162 1657 254 1691
<< labels >>
flabel locali s 990 689 1098 719 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 162 249 270 279 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 378 2053 486 2083 0 FreeSans 400 0 0 0 Q
port 4 nsew signal bidirectional
flabel locali s 378 1877 486 1907 0 FreeSans 400 0 0 0 QN
port 5 nsew signal bidirectional
flabel m3 s 774 0 874 2112 0 FreeSans 400 0 0 0 AVDD
port 6 nsew signal bidirectional
flabel m3 s 378 0 478 2112 0 FreeSans 400 0 0 0 AVSS
port 7 nsew signal bidirectional
flabel locali s 162 1657 270 1687 0 FreeSans 400 0 0 0 RN
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 2112
<< end >>
