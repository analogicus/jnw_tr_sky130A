magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 100 100
<< m2 >>
rect 0 0 100 100
<< v2 >>
rect 6 6 38 38
rect 6 62 38 94
rect 62 6 94 38
rect 62 62 94 94
<< m3 >>
rect 0 0 100 100
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 100 100
<< end >>
