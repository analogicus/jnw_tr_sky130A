magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1260 352
<< locali >>
rect 432 29 516 59
rect 516 29 828 59
rect 516 29 546 59
rect 432 293 516 323
rect 516 293 828 323
rect 516 293 546 323
rect 432 205 516 235
rect 516 205 828 235
rect 516 205 546 235
rect 201 73 231 191
rect 216 249 300 279
rect 300 29 432 59
rect 300 29 330 279
rect 1044 73 1128 103
rect 1044 249 1128 279
rect 1128 73 1158 279
rect 990 73 1098 103
rect 774 205 882 235
rect 378 293 486 323
<< poly >>
rect 162 79 1098 97
<< m3 >>
rect 828 117 918 155
rect 918 161 1044 199
rect 918 117 956 199
rect 774 0 874 352
rect 378 0 478 352
rect 774 0 874 352
rect 378 0 478 352
use JNWTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 630 176
use JNWTR_NCHDL MN1 
transform 1 0 0 0 1 88
box 0 88 630 264
use JNWTR_NCHDL MN2 
transform 1 0 0 0 1 176
box 0 176 630 352
use JNWTR_PCHDL MP0 
transform 1 0 630 0 1 0
box 630 0 1260 176
use JNWTR_PCHDL MP1_DMY 
transform 1 0 630 0 1 88
box 630 88 1260 264
use JNWTR_PCHDL MP2 
transform 1 0 630 0 1 176
box 630 176 1260 352
use JNWTR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 117
box 774 117 874 155
use JNWTR_cut_M1M4_2x1 xcut1 
transform 1 0 990 0 1 161
box 990 161 1090 199
use JNWTR_cut_M1M4_2x1 xcut2 
transform 1 0 774 0 1 117
box 774 117 874 155
use JNWTR_cut_M1M4_2x1 xcut3 
transform 1 0 378 0 1 117
box 378 117 478 155
use JNWTR_cut_M1M4_2x1 xcut4 
transform 1 0 378 0 1 117
box 378 117 478 155
<< labels >>
flabel locali s 990 73 1098 103 0 FreeSans 400 0 0 0 C
port 1 nsew signal bidirectional
flabel locali s 774 205 882 235 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 378 293 486 323 0 FreeSans 400 0 0 0 A
port 2 nsew signal bidirectional
flabel m3 s 774 0 874 352 0 FreeSans 400 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel m3 s 378 0 478 352 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 352
<< end >>
