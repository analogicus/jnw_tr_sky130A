magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1336 2118
<< locali >>
rect 8 8 1328 64
rect 64 8 1272 64
rect 8 8 1328 64
rect 64 2054 1272 2110
rect 8 2054 1328 2110
rect 8 64 64 2054
rect 8 8 64 2110
rect 1272 64 1328 2054
rect 1272 8 1328 2110
rect 8 8 1328 64
rect 740 1719 1028 1829
rect 308 1719 596 1829
<< ptapc >>
rect 88 16 128 56
rect 128 16 168 56
rect 168 16 208 56
rect 208 16 248 56
rect 248 16 288 56
rect 288 16 328 56
rect 328 16 368 56
rect 368 16 408 56
rect 408 16 448 56
rect 448 16 488 56
rect 488 16 528 56
rect 528 16 568 56
rect 568 16 608 56
rect 608 16 648 56
rect 648 16 688 56
rect 688 16 728 56
rect 728 16 768 56
rect 768 16 808 56
rect 808 16 848 56
rect 848 16 888 56
rect 888 16 928 56
rect 928 16 968 56
rect 968 16 1008 56
rect 1008 16 1048 56
rect 1048 16 1088 56
rect 1088 16 1128 56
rect 1128 16 1168 56
rect 1168 16 1208 56
rect 1208 16 1248 56
rect 88 2062 128 2102
rect 128 2062 168 2102
rect 168 2062 208 2102
rect 208 2062 248 2102
rect 248 2062 288 2102
rect 288 2062 328 2102
rect 328 2062 368 2102
rect 368 2062 408 2102
rect 408 2062 448 2102
rect 448 2062 488 2102
rect 488 2062 528 2102
rect 528 2062 568 2102
rect 568 2062 608 2102
rect 608 2062 648 2102
rect 648 2062 688 2102
rect 688 2062 728 2102
rect 728 2062 768 2102
rect 768 2062 808 2102
rect 808 2062 848 2102
rect 848 2062 888 2102
rect 888 2062 928 2102
rect 928 2062 968 2102
rect 968 2062 1008 2102
rect 1008 2062 1048 2102
rect 1048 2062 1088 2102
rect 1088 2062 1128 2102
rect 1128 2062 1168 2102
rect 1168 2062 1208 2102
rect 1208 2062 1248 2102
rect 16 79 56 119
rect 16 119 56 159
rect 16 159 56 199
rect 16 199 56 239
rect 16 239 56 279
rect 16 279 56 319
rect 16 319 56 359
rect 16 359 56 399
rect 16 399 56 439
rect 16 439 56 479
rect 16 479 56 519
rect 16 519 56 559
rect 16 559 56 599
rect 16 599 56 639
rect 16 639 56 679
rect 16 679 56 719
rect 16 719 56 759
rect 16 759 56 799
rect 16 799 56 839
rect 16 839 56 879
rect 16 879 56 919
rect 16 919 56 959
rect 16 959 56 999
rect 16 999 56 1039
rect 16 1039 56 1079
rect 16 1079 56 1119
rect 16 1119 56 1159
rect 16 1159 56 1199
rect 16 1199 56 1239
rect 16 1239 56 1279
rect 16 1279 56 1319
rect 16 1319 56 1359
rect 16 1359 56 1399
rect 16 1399 56 1439
rect 16 1439 56 1479
rect 16 1479 56 1519
rect 16 1519 56 1559
rect 16 1559 56 1599
rect 16 1599 56 1639
rect 16 1639 56 1679
rect 16 1679 56 1719
rect 16 1719 56 1759
rect 16 1759 56 1799
rect 16 1799 56 1839
rect 16 1839 56 1879
rect 16 1879 56 1919
rect 16 1919 56 1959
rect 16 1959 56 1999
rect 16 1999 56 2039
rect 1280 79 1320 119
rect 1280 119 1320 159
rect 1280 159 1320 199
rect 1280 199 1320 239
rect 1280 239 1320 279
rect 1280 279 1320 319
rect 1280 319 1320 359
rect 1280 359 1320 399
rect 1280 399 1320 439
rect 1280 439 1320 479
rect 1280 479 1320 519
rect 1280 519 1320 559
rect 1280 559 1320 599
rect 1280 599 1320 639
rect 1280 639 1320 679
rect 1280 679 1320 719
rect 1280 719 1320 759
rect 1280 759 1320 799
rect 1280 799 1320 839
rect 1280 839 1320 879
rect 1280 879 1320 919
rect 1280 919 1320 959
rect 1280 959 1320 999
rect 1280 999 1320 1039
rect 1280 1039 1320 1079
rect 1280 1079 1320 1119
rect 1280 1119 1320 1159
rect 1280 1159 1320 1199
rect 1280 1199 1320 1239
rect 1280 1239 1320 1279
rect 1280 1279 1320 1319
rect 1280 1319 1320 1359
rect 1280 1359 1320 1399
rect 1280 1399 1320 1439
rect 1280 1439 1320 1479
rect 1280 1479 1320 1519
rect 1280 1519 1320 1559
rect 1280 1559 1320 1599
rect 1280 1599 1320 1639
rect 1280 1639 1320 1679
rect 1280 1679 1320 1719
rect 1280 1719 1320 1759
rect 1280 1759 1320 1799
rect 1280 1799 1320 1839
rect 1280 1839 1320 1879
rect 1280 1879 1320 1919
rect 1280 1919 1320 1959
rect 1280 1959 1320 1999
rect 1280 1999 1320 2039
<< ptap >>
rect 0 0 1336 72
rect 0 2046 1336 2118
rect 0 0 72 2118
rect 1264 0 1336 2118
use JNWTR_RES2 XA1 
transform 1 0 344 0 1 344
box 344 344 992 1774
<< labels >>
flabel locali s 8 8 1328 64 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 740 1719 1028 1829 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel locali s 308 1719 596 1829 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1336 2118
<< end >>
