magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1944 1430
<< ppolyres >>
rect 180 -55 252 55
rect 396 -55 468 55
rect 612 -55 684 55
rect 828 -55 900 55
rect 1044 -55 1116 55
rect 1260 -55 1332 55
rect 1476 -55 1548 55
rect 1692 -55 1764 55
rect 180 55 252 165
rect 396 55 468 165
rect 612 55 684 165
rect 828 55 900 165
rect 1044 55 1116 165
rect 1260 55 1332 165
rect 1476 55 1548 165
rect 1692 55 1764 165
rect 180 165 252 275
rect 396 165 468 275
rect 612 165 684 275
rect 828 165 900 275
rect 1044 165 1116 275
rect 1260 165 1332 275
rect 1476 165 1548 275
rect 1692 165 1764 275
rect 180 275 252 385
rect 396 275 468 385
rect 612 275 684 385
rect 828 275 900 385
rect 1044 275 1116 385
rect 1260 275 1332 385
rect 1476 275 1548 385
rect 1692 275 1764 385
rect 180 385 252 495
rect 396 385 468 495
rect 612 385 684 495
rect 828 385 900 495
rect 1044 385 1116 495
rect 1260 385 1332 495
rect 1476 385 1548 495
rect 1692 385 1764 495
rect 180 495 252 605
rect 396 495 468 605
rect 612 495 684 605
rect 828 495 900 605
rect 1044 495 1116 605
rect 1260 495 1332 605
rect 1476 495 1548 605
rect 1692 495 1764 605
rect 180 605 252 715
rect 396 605 468 715
rect 612 605 684 715
rect 828 605 900 715
rect 1044 605 1116 715
rect 1260 605 1332 715
rect 1476 605 1548 715
rect 1692 605 1764 715
rect 180 715 252 825
rect 396 715 468 825
rect 612 715 684 825
rect 828 715 900 825
rect 1044 715 1116 825
rect 1260 715 1332 825
rect 1476 715 1548 825
rect 1692 715 1764 825
rect 180 825 252 935
rect 396 825 468 935
rect 612 825 684 935
rect 828 825 900 935
rect 1044 825 1116 935
rect 1260 825 1332 935
rect 1476 825 1548 935
rect 1692 825 1764 935
rect 180 935 252 1045
rect 396 935 468 1045
rect 612 935 684 1045
rect 828 935 900 1045
rect 1044 935 1116 1045
rect 1260 935 1332 1045
rect 1476 935 1548 1045
rect 1692 935 1764 1045
rect 180 1045 252 1155
rect 396 1045 468 1155
rect 612 1045 684 1155
rect 828 1045 900 1155
rect 1044 1045 1116 1155
rect 1260 1045 1332 1155
rect 1476 1045 1548 1155
rect 1692 1045 1764 1155
rect 180 1155 252 1265
rect 396 1155 468 1265
rect 612 1155 684 1265
rect 828 1155 900 1265
rect 1044 1155 1116 1265
rect 1260 1155 1332 1265
rect 1476 1155 1548 1265
rect 1692 1155 1764 1265
<< poly >>
rect -36 -55 36 55
rect 1908 -55 1980 55
rect -36 55 36 165
rect 1908 55 1980 165
rect -36 165 36 275
rect 1908 165 1980 275
rect -36 275 36 385
rect 1908 275 1980 385
rect -36 385 36 495
rect 1908 385 1980 495
rect -36 495 36 605
rect 1908 495 1980 605
rect -36 605 36 715
rect 1908 605 1980 715
rect -36 715 36 825
rect 1908 715 1980 825
rect -36 825 36 935
rect 1908 825 1980 935
rect -36 935 36 1045
rect 1908 935 1980 1045
rect -36 1045 36 1155
rect 1908 1045 1980 1155
rect -36 1155 36 1265
rect 1908 1155 1980 1265
<< xpolycontact >>
rect 180 -55 252 55
rect 396 -55 468 55
rect 612 -55 684 55
rect 828 -55 900 55
rect 1044 -55 1116 55
rect 1260 -55 1332 55
rect 1476 -55 1548 55
rect 1692 -55 1764 55
rect 180 55 252 165
rect 396 55 468 165
rect 612 55 684 165
rect 828 55 900 165
rect 1044 55 1116 165
rect 1260 55 1332 165
rect 1476 55 1548 165
rect 1692 55 1764 165
rect 180 1045 252 1155
rect 396 1045 468 1155
rect 612 1045 684 1155
rect 828 1045 900 1155
rect 1044 1045 1116 1155
rect 1260 1045 1332 1155
rect 1476 1045 1548 1155
rect 1692 1045 1764 1155
rect 180 1155 252 1265
rect 396 1155 468 1265
rect 612 1155 684 1265
rect 828 1155 900 1265
rect 1044 1155 1116 1265
rect 1260 1155 1332 1265
rect 1476 1155 1548 1265
rect 1692 1155 1764 1265
<< locali >>
rect 180 -55 468 55
rect 612 -55 900 55
rect 1044 -55 1332 55
rect 1476 -55 1764 55
rect 180 55 468 165
rect 612 55 900 165
rect 1044 55 1332 165
rect 1476 55 1764 165
rect 180 1045 252 1155
rect 396 1045 468 1155
rect 612 1045 684 1155
rect 828 1045 900 1155
rect 1044 1045 1116 1155
rect 1260 1045 1332 1155
rect 1476 1045 1548 1155
rect 1692 1045 1764 1155
rect 180 1155 252 1265
rect 396 1155 468 1265
rect 612 1155 684 1265
rect 828 1155 900 1265
rect 1044 1155 1116 1265
rect 1260 1155 1332 1265
rect 1476 1155 1548 1265
rect 1692 1155 1764 1265
rect 180 1265 252 1375
rect 396 1265 468 1375
rect 612 1265 684 1375
rect 828 1265 900 1375
rect 1044 1265 1116 1375
rect 1260 1265 1332 1375
rect 1476 1265 1548 1375
rect 1692 1265 1764 1375
rect -36 1375 252 1485
rect -36 1375 252 1485
rect 396 1375 684 1485
rect 828 1375 1116 1485
rect 1260 1375 1548 1485
rect 1692 1375 1980 1485
rect 1692 1375 1980 1485
<< pwell >>
rect -36 -55 1980 1485
<< labels >>
flabel locali s -36 1375 252 1485 0 FreeSans 400 0 0 0 N
port 1 nsew signal bidirectional
flabel locali s 1692 1375 1980 1485 0 FreeSans 400 0 0 0 P
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1944 1430
<< end >>
