magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1260 528
<< locali >>
rect 417 293 447 411
rect 813 117 843 235
rect 432 205 516 235
rect 516 469 828 499
rect 516 205 546 499
rect 102 425 216 455
rect 102 147 408 177
rect 102 147 132 455
rect 378 117 432 147
rect 432 117 582 147
rect 582 293 828 323
rect 582 117 612 323
rect 162 73 270 103
rect 162 249 270 279
rect 378 205 486 235
<< poly >>
rect 162 79 1098 97
rect 162 255 1098 273
rect 162 431 1098 449
<< m3 >>
rect 774 0 874 528
rect 378 0 478 528
rect 774 0 874 528
rect 378 0 478 528
use JNWTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 630 176
use JNWTR_NCHDL MN2 
transform 1 0 0 0 1 176
box 0 176 630 352
use JNWTR_NCHDL MN1 
transform 1 0 0 0 1 352
box 0 352 630 528
use JNWTR_PCHDL MP1 
transform 1 0 630 0 1 0
box 630 0 1260 176
use JNWTR_PCHDL MP0 
transform 1 0 630 0 1 176
box 630 176 1260 352
use JNWTR_PCHDL MP2 
transform 1 0 630 0 1 352
box 630 352 1260 528
use JNWTR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 29
box 774 29 874 67
use JNWTR_cut_M1M4_2x1 xcut1 
transform 1 0 774 0 1 381
box 774 381 874 419
use JNWTR_cut_M1M4_2x1 xcut2 
transform 1 0 378 0 1 29
box 378 29 478 67
use JNWTR_cut_M1M4_2x1 xcut3 
transform 1 0 378 0 1 469
box 378 469 478 507
<< labels >>
flabel locali s 162 73 270 103 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
flabel locali s 162 249 270 279 0 FreeSans 400 0 0 0 CK
port 2 nsew signal bidirectional
flabel locali s 378 205 486 235 0 FreeSans 400 0 0 0 Q
port 3 nsew signal bidirectional
flabel m3 s 774 0 874 528 0 FreeSans 400 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel m3 s 378 0 478 528 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 528
<< end >>
