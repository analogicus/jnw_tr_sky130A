magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 1836 1320
<< ppolyres >>
rect 90 -60 126 60
rect 198 -60 234 60
rect 306 -60 342 60
rect 414 -60 450 60
rect 522 -60 558 60
rect 630 -60 666 60
rect 738 -60 774 60
rect 846 -60 882 60
rect 954 -60 990 60
rect 1062 -60 1098 60
rect 1170 -60 1206 60
rect 1278 -60 1314 60
rect 1386 -60 1422 60
rect 1494 -60 1530 60
rect 1602 -60 1638 60
rect 1710 -60 1746 60
rect 90 60 126 180
rect 198 60 234 180
rect 306 60 342 180
rect 414 60 450 180
rect 522 60 558 180
rect 630 60 666 180
rect 738 60 774 180
rect 846 60 882 180
rect 954 60 990 180
rect 1062 60 1098 180
rect 1170 60 1206 180
rect 1278 60 1314 180
rect 1386 60 1422 180
rect 1494 60 1530 180
rect 1602 60 1638 180
rect 1710 60 1746 180
rect 90 180 126 300
rect 198 180 234 300
rect 306 180 342 300
rect 414 180 450 300
rect 522 180 558 300
rect 630 180 666 300
rect 738 180 774 300
rect 846 180 882 300
rect 954 180 990 300
rect 1062 180 1098 300
rect 1170 180 1206 300
rect 1278 180 1314 300
rect 1386 180 1422 300
rect 1494 180 1530 300
rect 1602 180 1638 300
rect 1710 180 1746 300
rect 90 300 126 420
rect 198 300 234 420
rect 306 300 342 420
rect 414 300 450 420
rect 522 300 558 420
rect 630 300 666 420
rect 738 300 774 420
rect 846 300 882 420
rect 954 300 990 420
rect 1062 300 1098 420
rect 1170 300 1206 420
rect 1278 300 1314 420
rect 1386 300 1422 420
rect 1494 300 1530 420
rect 1602 300 1638 420
rect 1710 300 1746 420
rect 90 420 126 540
rect 198 420 234 540
rect 306 420 342 540
rect 414 420 450 540
rect 522 420 558 540
rect 630 420 666 540
rect 738 420 774 540
rect 846 420 882 540
rect 954 420 990 540
rect 1062 420 1098 540
rect 1170 420 1206 540
rect 1278 420 1314 540
rect 1386 420 1422 540
rect 1494 420 1530 540
rect 1602 420 1638 540
rect 1710 420 1746 540
rect 90 540 126 660
rect 198 540 234 660
rect 306 540 342 660
rect 414 540 450 660
rect 522 540 558 660
rect 630 540 666 660
rect 738 540 774 660
rect 846 540 882 660
rect 954 540 990 660
rect 1062 540 1098 660
rect 1170 540 1206 660
rect 1278 540 1314 660
rect 1386 540 1422 660
rect 1494 540 1530 660
rect 1602 540 1638 660
rect 1710 540 1746 660
rect 90 660 126 780
rect 198 660 234 780
rect 306 660 342 780
rect 414 660 450 780
rect 522 660 558 780
rect 630 660 666 780
rect 738 660 774 780
rect 846 660 882 780
rect 954 660 990 780
rect 1062 660 1098 780
rect 1170 660 1206 780
rect 1278 660 1314 780
rect 1386 660 1422 780
rect 1494 660 1530 780
rect 1602 660 1638 780
rect 1710 660 1746 780
rect 90 780 126 900
rect 198 780 234 900
rect 306 780 342 900
rect 414 780 450 900
rect 522 780 558 900
rect 630 780 666 900
rect 738 780 774 900
rect 846 780 882 900
rect 954 780 990 900
rect 1062 780 1098 900
rect 1170 780 1206 900
rect 1278 780 1314 900
rect 1386 780 1422 900
rect 1494 780 1530 900
rect 1602 780 1638 900
rect 1710 780 1746 900
rect 90 900 126 1020
rect 198 900 234 1020
rect 306 900 342 1020
rect 414 900 450 1020
rect 522 900 558 1020
rect 630 900 666 1020
rect 738 900 774 1020
rect 846 900 882 1020
rect 954 900 990 1020
rect 1062 900 1098 1020
rect 1170 900 1206 1020
rect 1278 900 1314 1020
rect 1386 900 1422 1020
rect 1494 900 1530 1020
rect 1602 900 1638 1020
rect 1710 900 1746 1020
rect 90 1020 126 1140
rect 198 1020 234 1140
rect 306 1020 342 1140
rect 414 1020 450 1140
rect 522 1020 558 1140
rect 630 1020 666 1140
rect 738 1020 774 1140
rect 846 1020 882 1140
rect 954 1020 990 1140
rect 1062 1020 1098 1140
rect 1170 1020 1206 1140
rect 1278 1020 1314 1140
rect 1386 1020 1422 1140
rect 1494 1020 1530 1140
rect 1602 1020 1638 1140
rect 1710 1020 1746 1140
<< poly >>
rect -18 -60 18 60
rect 1818 -60 1854 60
rect -18 60 18 180
rect 1818 60 1854 180
rect -18 180 18 300
rect 1818 180 1854 300
rect -18 300 18 420
rect 1818 300 1854 420
rect -18 420 18 540
rect 1818 420 1854 540
rect -18 540 18 660
rect 1818 540 1854 660
rect -18 660 18 780
rect 1818 660 1854 780
rect -18 780 18 900
rect 1818 780 1854 900
rect -18 900 18 1020
rect 1818 900 1854 1020
rect -18 1020 18 1140
rect 1818 1020 1854 1140
<< xpolycontact >>
rect 90 -60 126 60
rect 198 -60 234 60
rect 306 -60 342 60
rect 414 -60 450 60
rect 522 -60 558 60
rect 630 -60 666 60
rect 738 -60 774 60
rect 846 -60 882 60
rect 954 -60 990 60
rect 1062 -60 1098 60
rect 1170 -60 1206 60
rect 1278 -60 1314 60
rect 1386 -60 1422 60
rect 1494 -60 1530 60
rect 1602 -60 1638 60
rect 1710 -60 1746 60
rect 90 60 126 180
rect 198 60 234 180
rect 306 60 342 180
rect 414 60 450 180
rect 522 60 558 180
rect 630 60 666 180
rect 738 60 774 180
rect 846 60 882 180
rect 954 60 990 180
rect 1062 60 1098 180
rect 1170 60 1206 180
rect 1278 60 1314 180
rect 1386 60 1422 180
rect 1494 60 1530 180
rect 1602 60 1638 180
rect 1710 60 1746 180
rect 90 900 126 1020
rect 198 900 234 1020
rect 306 900 342 1020
rect 414 900 450 1020
rect 522 900 558 1020
rect 630 900 666 1020
rect 738 900 774 1020
rect 846 900 882 1020
rect 954 900 990 1020
rect 1062 900 1098 1020
rect 1170 900 1206 1020
rect 1278 900 1314 1020
rect 1386 900 1422 1020
rect 1494 900 1530 1020
rect 1602 900 1638 1020
rect 1710 900 1746 1020
rect 90 1020 126 1140
rect 198 1020 234 1140
rect 306 1020 342 1140
rect 414 1020 450 1140
rect 522 1020 558 1140
rect 630 1020 666 1140
rect 738 1020 774 1140
rect 846 1020 882 1140
rect 954 1020 990 1140
rect 1062 1020 1098 1140
rect 1170 1020 1206 1140
rect 1278 1020 1314 1140
rect 1386 1020 1422 1140
rect 1494 1020 1530 1140
rect 1602 1020 1638 1140
rect 1710 1020 1746 1140
<< locali >>
rect 90 -60 234 60
rect 306 -60 450 60
rect 522 -60 666 60
rect 738 -60 882 60
rect 954 -60 1098 60
rect 1170 -60 1314 60
rect 1386 -60 1530 60
rect 1602 -60 1746 60
rect 90 60 234 180
rect 306 60 450 180
rect 522 60 666 180
rect 738 60 882 180
rect 954 60 1098 180
rect 1170 60 1314 180
rect 1386 60 1530 180
rect 1602 60 1746 180
rect 90 900 126 1020
rect 198 900 234 1020
rect 306 900 342 1020
rect 414 900 450 1020
rect 522 900 558 1020
rect 630 900 666 1020
rect 738 900 774 1020
rect 846 900 882 1020
rect 954 900 990 1020
rect 1062 900 1098 1020
rect 1170 900 1206 1020
rect 1278 900 1314 1020
rect 1386 900 1422 1020
rect 1494 900 1530 1020
rect 1602 900 1638 1020
rect 1710 900 1746 1020
rect 90 1020 126 1140
rect 198 1020 234 1140
rect 306 1020 342 1140
rect 414 1020 450 1140
rect 522 1020 558 1140
rect 630 1020 666 1140
rect 738 1020 774 1140
rect 846 1020 882 1140
rect 954 1020 990 1140
rect 1062 1020 1098 1140
rect 1170 1020 1206 1140
rect 1278 1020 1314 1140
rect 1386 1020 1422 1140
rect 1494 1020 1530 1140
rect 1602 1020 1638 1140
rect 1710 1020 1746 1140
rect 90 1140 126 1260
rect 198 1140 234 1260
rect 306 1140 342 1260
rect 414 1140 450 1260
rect 522 1140 558 1260
rect 630 1140 666 1260
rect 738 1140 774 1260
rect 846 1140 882 1260
rect 954 1140 990 1260
rect 1062 1140 1098 1260
rect 1170 1140 1206 1260
rect 1278 1140 1314 1260
rect 1386 1140 1422 1260
rect 1494 1140 1530 1260
rect 1602 1140 1638 1260
rect 1710 1140 1746 1260
rect -18 1260 126 1380
rect -18 1260 126 1380
rect 198 1260 342 1380
rect 414 1260 558 1380
rect 630 1260 774 1380
rect 846 1260 990 1380
rect 1062 1260 1206 1380
rect 1278 1260 1422 1380
rect 1494 1260 1638 1380
rect 1710 1260 1854 1380
rect 1710 1260 1854 1380
<< pwell >>
rect -18 -60 1854 1380
<< labels >>
flabel locali s -18 1260 126 1380 0 FreeSans 400 0 0 0 N
port 1 nsew signal bidirectional
flabel locali s 1710 1260 1854 1380 0 FreeSans 400 0 0 0 P
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1836 1320
<< end >>
