magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1260 176
<< locali >>
rect 216 73 300 103
rect 300 117 432 147
rect 300 73 330 147
rect 774 117 882 147
<< poly >>
rect 162 79 1098 97
<< m3 >>
rect 774 0 874 176
rect 378 0 478 176
rect 774 0 874 176
rect 378 0 478 176
use JNWTR_NCHDL MN0 
transform 1 0 0 0 1 0
box 0 0 630 176
use JNWTR_PCHDL MP0 
transform 1 0 630 0 1 0
box 630 0 1260 176
use JNWTR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 29
box 774 29 874 67
use JNWTR_cut_M1M4_2x1 xcut1 
transform 1 0 378 0 1 29
box 378 29 478 67
<< labels >>
flabel locali s 774 117 882 147 0 FreeSans 400 0 0 0 Y
port 1 nsew signal bidirectional
flabel m3 s 774 0 874 176 0 FreeSans 400 0 0 0 AVDD
port 2 nsew signal bidirectional
flabel m3 s 378 0 478 176 0 FreeSans 400 0 0 0 AVSS
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 176
<< end >>
