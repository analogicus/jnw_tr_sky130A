magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1260 440
<< locali >>
rect 216 337 300 367
rect 300 205 432 235
rect 300 205 330 367
rect 162 73 270 103
rect 162 161 270 191
rect 378 381 486 411
<< m3 >>
rect 774 0 874 440
rect 378 0 478 440
rect 774 0 874 440
rect 378 0 478 440
use JNWTR_NDX1_CV XA1 
transform 1 0 0 0 1 0
box 0 0 1260 264
use JNWTR_IVX1_CV XA2 
transform 1 0 0 0 1 264
box 0 264 1260 440
<< labels >>
flabel locali s 162 73 270 103 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 162 161 270 191 0 FreeSans 400 0 0 0 B
port 2 nsew signal bidirectional
flabel locali s 378 381 486 411 0 FreeSans 400 0 0 0 Y
port 3 nsew signal bidirectional
flabel m3 s 774 0 874 440 0 FreeSans 400 0 0 0 AVDD
port 4 nsew signal bidirectional
flabel m3 s 378 0 478 440 0 FreeSans 400 0 0 0 AVSS
port 5 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 440
<< end >>
