magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 88 34
<< locali >>
rect 0 0 84 32
<< viali >>
rect 6 3 32 29
rect 52 3 78 29
<< m1 >>
rect 0 0 88 34
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 88 34
<< end >>
