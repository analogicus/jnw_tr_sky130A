magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1260 880
<< locali >>
rect 432 117 516 147
rect 432 205 516 235
rect 432 381 516 411
rect 432 557 516 587
rect 516 117 546 587
rect 714 117 828 147
rect 714 205 828 235
rect 714 469 828 499
rect 714 645 828 675
rect 714 117 744 675
rect 201 73 231 279
rect 1044 425 1128 455
rect 852 323 1128 353
rect 1068 631 1128 661
rect 1068 807 1128 837
rect 1128 323 1158 837
rect 828 293 882 323
rect 1044 601 1098 631
rect 1044 777 1098 807
rect 102 425 216 455
rect 102 323 408 353
rect 102 631 192 661
rect 102 807 192 837
rect 102 323 132 837
rect 378 293 432 323
rect 162 601 216 631
rect 162 777 216 807
rect 318 469 432 499
rect 318 645 432 675
rect 318 469 348 675
rect 432 821 516 851
rect 516 821 828 851
rect 516 821 546 851
rect 432 645 516 675
rect 516 733 828 763
rect 516 645 546 763
rect 828 381 912 411
rect 828 557 912 587
rect 912 381 942 587
rect 162 73 270 103
rect 378 821 486 851
<< m1 >>
rect 432 733 516 763
rect 516 557 828 587
rect 516 557 546 763
rect 432 293 516 323
rect 516 293 828 323
rect 516 293 546 323
<< poly >>
rect 162 79 1098 97
rect 162 255 1098 273
<< m3 >>
rect 774 0 874 880
rect 378 0 478 880
rect 774 0 874 880
rect 378 0 478 880
use JNWTR_NCHDL XA2 
transform 1 0 0 0 1 0
box 0 0 630 176
use JNWTR_NCHDL XA3 
transform 1 0 0 0 1 176
box 0 176 630 352
use JNWTR_NCHDL XA4a 
transform 1 0 0 0 1 352
box 0 352 630 528
use JNWTR_NCHDL XA4b 
transform 1 0 0 0 1 528
box 0 528 630 704
use JNWTR_NCHDL XA5 
transform 1 0 0 0 1 704
box 0 704 630 880
use JNWTR_PCHDL XB0 
transform 1 0 630 0 1 0
box 630 0 1260 176
use JNWTR_PCHDL XB1 
transform 1 0 630 0 1 176
box 630 176 1260 352
use JNWTR_PCHDL XB3a 
transform 1 0 630 0 1 352
box 630 352 1260 528
use JNWTR_PCHDL XB3b 
transform 1 0 630 0 1 528
box 630 528 1260 704
use JNWTR_PCHDL XB4 
transform 1 0 630 0 1 704
box 630 704 1260 880
use JNWTR_cut_M1M2_2x1 xcut0 
transform 1 0 378 0 1 733
box 378 733 470 767
use JNWTR_cut_M1M2_2x1 xcut1 
transform 1 0 774 0 1 557
box 774 557 866 591
use JNWTR_cut_M1M2_2x1 xcut2 
transform 1 0 378 0 1 293
box 378 293 470 327
use JNWTR_cut_M1M2_2x1 xcut3 
transform 1 0 774 0 1 293
box 774 293 866 327
use JNWTR_cut_M1M4_2x1 xcut4 
transform 1 0 774 0 1 29
box 774 29 874 67
use JNWTR_cut_M1M4_2x1 xcut5 
transform 1 0 774 0 1 733
box 774 733 874 771
use JNWTR_cut_M1M4_2x1 xcut6 
transform 1 0 378 0 1 29
box 378 29 478 67
use JNWTR_cut_M1M4_2x1 xcut7 
transform 1 0 378 0 1 733
box 378 733 478 771
<< labels >>
flabel locali s 162 73 270 103 0 FreeSans 400 0 0 0 A
port 1 nsew signal bidirectional
flabel locali s 378 821 486 851 0 FreeSans 400 0 0 0 Y
port 2 nsew signal bidirectional
flabel m3 s 774 0 874 880 0 FreeSans 400 0 0 0 AVDD
port 3 nsew signal bidirectional
flabel m3 s 378 0 478 880 0 FreeSans 400 0 0 0 AVSS
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 880
<< end >>
