magic
tech sky130A
magscale 1 1
timestamp 1723932000
<< checkpaint >>
rect 0 0 1372 1720
<< locali >>
rect 8 8 1364 64
rect 64 8 1308 64
rect 8 8 1364 64
rect 64 1656 1308 1712
rect 8 1656 1364 1712
rect 8 64 64 1656
rect 8 8 64 1712
rect 1308 64 1364 1656
rect 1308 8 1364 1712
rect 8 8 1364 64
rect 1046 1460 1190 1580
rect 182 1460 326 1580
<< ptapc >>
rect 86 16 126 56
rect 126 16 166 56
rect 166 16 206 56
rect 206 16 246 56
rect 246 16 286 56
rect 286 16 326 56
rect 326 16 366 56
rect 366 16 406 56
rect 406 16 446 56
rect 446 16 486 56
rect 486 16 526 56
rect 526 16 566 56
rect 566 16 606 56
rect 606 16 646 56
rect 646 16 686 56
rect 686 16 726 56
rect 726 16 766 56
rect 766 16 806 56
rect 806 16 846 56
rect 846 16 886 56
rect 886 16 926 56
rect 926 16 966 56
rect 966 16 1006 56
rect 1006 16 1046 56
rect 1046 16 1086 56
rect 1086 16 1126 56
rect 1126 16 1166 56
rect 1166 16 1206 56
rect 1206 16 1246 56
rect 1246 16 1286 56
rect 86 1664 126 1704
rect 126 1664 166 1704
rect 166 1664 206 1704
rect 206 1664 246 1704
rect 246 1664 286 1704
rect 286 1664 326 1704
rect 326 1664 366 1704
rect 366 1664 406 1704
rect 406 1664 446 1704
rect 446 1664 486 1704
rect 486 1664 526 1704
rect 526 1664 566 1704
rect 566 1664 606 1704
rect 606 1664 646 1704
rect 646 1664 686 1704
rect 686 1664 726 1704
rect 726 1664 766 1704
rect 766 1664 806 1704
rect 806 1664 846 1704
rect 846 1664 886 1704
rect 886 1664 926 1704
rect 926 1664 966 1704
rect 966 1664 1006 1704
rect 1006 1664 1046 1704
rect 1046 1664 1086 1704
rect 1086 1664 1126 1704
rect 1126 1664 1166 1704
rect 1166 1664 1206 1704
rect 1206 1664 1246 1704
rect 1246 1664 1286 1704
rect 16 80 56 120
rect 16 120 56 160
rect 16 160 56 200
rect 16 200 56 240
rect 16 240 56 280
rect 16 280 56 320
rect 16 320 56 360
rect 16 360 56 400
rect 16 400 56 440
rect 16 440 56 480
rect 16 480 56 520
rect 16 520 56 560
rect 16 560 56 600
rect 16 600 56 640
rect 16 640 56 680
rect 16 680 56 720
rect 16 720 56 760
rect 16 760 56 800
rect 16 800 56 840
rect 16 840 56 880
rect 16 880 56 920
rect 16 920 56 960
rect 16 960 56 1000
rect 16 1000 56 1040
rect 16 1040 56 1080
rect 16 1080 56 1120
rect 16 1120 56 1160
rect 16 1160 56 1200
rect 16 1200 56 1240
rect 16 1240 56 1280
rect 16 1280 56 1320
rect 16 1320 56 1360
rect 16 1360 56 1400
rect 16 1400 56 1440
rect 16 1440 56 1480
rect 16 1480 56 1520
rect 16 1520 56 1560
rect 16 1560 56 1600
rect 16 1600 56 1640
rect 1316 80 1356 120
rect 1316 120 1356 160
rect 1316 160 1356 200
rect 1316 200 1356 240
rect 1316 240 1356 280
rect 1316 280 1356 320
rect 1316 320 1356 360
rect 1316 360 1356 400
rect 1316 400 1356 440
rect 1316 440 1356 480
rect 1316 480 1356 520
rect 1316 520 1356 560
rect 1316 560 1356 600
rect 1316 600 1356 640
rect 1316 640 1356 680
rect 1316 680 1356 720
rect 1316 720 1356 760
rect 1316 760 1356 800
rect 1316 800 1356 840
rect 1316 840 1356 880
rect 1316 880 1356 920
rect 1316 920 1356 960
rect 1316 960 1356 1000
rect 1316 1000 1356 1040
rect 1316 1040 1356 1080
rect 1316 1080 1356 1120
rect 1316 1120 1356 1160
rect 1316 1160 1356 1200
rect 1316 1200 1356 1240
rect 1316 1240 1356 1280
rect 1316 1280 1356 1320
rect 1316 1320 1356 1360
rect 1316 1360 1356 1400
rect 1316 1400 1356 1440
rect 1316 1440 1356 1480
rect 1316 1480 1356 1520
rect 1316 1520 1356 1560
rect 1316 1560 1356 1600
rect 1316 1600 1356 1640
<< ptap >>
rect 0 0 1372 72
rect 0 1648 1372 1720
rect 0 0 72 1720
rect 1300 0 1372 1720
use JNWTR_RES8 XA1 
transform 1 0 200 0 1 200
box 200 200 1172 1520
<< labels >>
flabel locali s 8 8 1364 64 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 1046 1460 1190 1580 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel locali s 182 1460 326 1580 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1372 1720
<< end >>
