magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 630 176
<< pdiff >>
rect 144 22 252 66
rect 144 66 252 110
rect 144 110 252 154
<< ntap >>
rect 576 -22 684 22
rect 576 22 684 66
rect 576 66 684 110
rect 576 110 684 154
rect 576 154 684 198
<< poly >>
rect 108 -9 468 9
rect 108 79 468 97
rect 108 167 468 185
rect 360 66 468 110
<< locali >>
rect 360 73 468 103
rect 576 -22 684 22
rect 144 29 252 59
rect 144 29 252 59
rect 576 22 684 66
rect 360 73 468 103
rect 576 66 684 110
rect 576 66 684 110
rect 144 117 252 147
rect 144 117 252 147
rect 576 110 684 154
rect 576 154 684 198
<< pcontact >>
rect 372 77 396 88
rect 372 88 396 99
rect 396 77 432 88
rect 396 88 432 99
rect 432 77 456 88
rect 432 88 456 99
<< ntapc >>
rect 612 22 648 66
rect 612 110 648 154
<< pdcontact >>
rect 156 33 180 44
rect 156 44 180 55
rect 180 33 216 44
rect 180 44 216 55
rect 216 33 240 44
rect 216 44 240 55
rect 156 121 180 132
rect 156 132 180 143
rect 180 121 216 132
rect 180 132 216 143
rect 216 121 240 132
rect 216 132 240 143
<< nwell >>
rect 0 -66 720 242
<< labels >>
flabel locali s 360 73 468 103 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel locali s 144 29 252 59 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel locali s 576 66 684 110 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel locali s 144 117 252 147 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 630 176
<< end >>
