magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 1260 176
<< locali >>
rect -54 73 270 103
rect 216 73 300 103
rect 300 29 432 59
rect 300 29 330 103
rect 216 73 300 103
rect 300 117 432 147
rect 300 73 330 147
rect 828 29 912 59
rect 912 73 1044 103
rect 912 29 942 103
rect 828 117 912 147
rect 912 73 1044 103
rect 912 73 942 147
rect 990 73 1314 103
<< m3 >>
rect 774 0 874 176
rect 378 0 478 176
rect 774 0 874 176
rect 378 0 478 176
use JNWTR_NCHDL MN1 
transform 1 0 0 0 1 0
box 0 0 630 176
use JNWTR_PCHDL MP1 
transform 1 0 630 0 1 0
box 630 0 1260 176
use JNWTR_cut_M1M4_2x1 xcut0 
transform 1 0 774 0 1 117
box 774 117 874 155
use JNWTR_cut_M1M4_2x1 xcut1 
transform 1 0 774 0 1 29
box 774 29 874 67
use JNWTR_cut_M1M4_2x1 xcut2 
transform 1 0 378 0 1 117
box 378 117 478 155
use JNWTR_cut_M1M4_2x1 xcut3 
transform 1 0 378 0 1 29
box 378 29 478 67
<< labels >>
flabel m3 s 774 0 874 176 0 FreeSans 400 0 0 0 AVDD
port 1 nsew signal bidirectional
flabel m3 s 378 0 478 176 0 FreeSans 400 0 0 0 AVSS
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1260 176
<< end >>
