magic
tech sky130A
magscale 1 1
timestamp 1723845600
<< checkpaint >>
rect 0 0 4360 2118
<< locali >>
rect 8 8 4352 64
rect 64 8 4296 64
rect 8 8 4352 64
rect 64 2054 4296 2110
rect 8 2054 4352 2110
rect 8 64 64 2054
rect 8 8 64 2110
rect 4296 64 4352 2054
rect 4296 8 4352 2110
rect 8 8 4352 64
rect 3764 1719 4052 1829
rect 308 1719 596 1829
<< ptapc >>
rect 80 16 120 56
rect 120 16 160 56
rect 160 16 200 56
rect 200 16 240 56
rect 240 16 280 56
rect 280 16 320 56
rect 320 16 360 56
rect 360 16 400 56
rect 400 16 440 56
rect 440 16 480 56
rect 480 16 520 56
rect 520 16 560 56
rect 560 16 600 56
rect 600 16 640 56
rect 640 16 680 56
rect 680 16 720 56
rect 720 16 760 56
rect 760 16 800 56
rect 800 16 840 56
rect 840 16 880 56
rect 880 16 920 56
rect 920 16 960 56
rect 960 16 1000 56
rect 1000 16 1040 56
rect 1040 16 1080 56
rect 1080 16 1120 56
rect 1120 16 1160 56
rect 1160 16 1200 56
rect 1200 16 1240 56
rect 1240 16 1280 56
rect 1280 16 1320 56
rect 1320 16 1360 56
rect 1360 16 1400 56
rect 1400 16 1440 56
rect 1440 16 1480 56
rect 1480 16 1520 56
rect 1520 16 1560 56
rect 1560 16 1600 56
rect 1600 16 1640 56
rect 1640 16 1680 56
rect 1680 16 1720 56
rect 1720 16 1760 56
rect 1760 16 1800 56
rect 1800 16 1840 56
rect 1840 16 1880 56
rect 1880 16 1920 56
rect 1920 16 1960 56
rect 1960 16 2000 56
rect 2000 16 2040 56
rect 2040 16 2080 56
rect 2080 16 2120 56
rect 2120 16 2160 56
rect 2160 16 2200 56
rect 2200 16 2240 56
rect 2240 16 2280 56
rect 2280 16 2320 56
rect 2320 16 2360 56
rect 2360 16 2400 56
rect 2400 16 2440 56
rect 2440 16 2480 56
rect 2480 16 2520 56
rect 2520 16 2560 56
rect 2560 16 2600 56
rect 2600 16 2640 56
rect 2640 16 2680 56
rect 2680 16 2720 56
rect 2720 16 2760 56
rect 2760 16 2800 56
rect 2800 16 2840 56
rect 2840 16 2880 56
rect 2880 16 2920 56
rect 2920 16 2960 56
rect 2960 16 3000 56
rect 3000 16 3040 56
rect 3040 16 3080 56
rect 3080 16 3120 56
rect 3120 16 3160 56
rect 3160 16 3200 56
rect 3200 16 3240 56
rect 3240 16 3280 56
rect 3280 16 3320 56
rect 3320 16 3360 56
rect 3360 16 3400 56
rect 3400 16 3440 56
rect 3440 16 3480 56
rect 3480 16 3520 56
rect 3520 16 3560 56
rect 3560 16 3600 56
rect 3600 16 3640 56
rect 3640 16 3680 56
rect 3680 16 3720 56
rect 3720 16 3760 56
rect 3760 16 3800 56
rect 3800 16 3840 56
rect 3840 16 3880 56
rect 3880 16 3920 56
rect 3920 16 3960 56
rect 3960 16 4000 56
rect 4000 16 4040 56
rect 4040 16 4080 56
rect 4080 16 4120 56
rect 4120 16 4160 56
rect 4160 16 4200 56
rect 4200 16 4240 56
rect 4240 16 4280 56
rect 80 2062 120 2102
rect 120 2062 160 2102
rect 160 2062 200 2102
rect 200 2062 240 2102
rect 240 2062 280 2102
rect 280 2062 320 2102
rect 320 2062 360 2102
rect 360 2062 400 2102
rect 400 2062 440 2102
rect 440 2062 480 2102
rect 480 2062 520 2102
rect 520 2062 560 2102
rect 560 2062 600 2102
rect 600 2062 640 2102
rect 640 2062 680 2102
rect 680 2062 720 2102
rect 720 2062 760 2102
rect 760 2062 800 2102
rect 800 2062 840 2102
rect 840 2062 880 2102
rect 880 2062 920 2102
rect 920 2062 960 2102
rect 960 2062 1000 2102
rect 1000 2062 1040 2102
rect 1040 2062 1080 2102
rect 1080 2062 1120 2102
rect 1120 2062 1160 2102
rect 1160 2062 1200 2102
rect 1200 2062 1240 2102
rect 1240 2062 1280 2102
rect 1280 2062 1320 2102
rect 1320 2062 1360 2102
rect 1360 2062 1400 2102
rect 1400 2062 1440 2102
rect 1440 2062 1480 2102
rect 1480 2062 1520 2102
rect 1520 2062 1560 2102
rect 1560 2062 1600 2102
rect 1600 2062 1640 2102
rect 1640 2062 1680 2102
rect 1680 2062 1720 2102
rect 1720 2062 1760 2102
rect 1760 2062 1800 2102
rect 1800 2062 1840 2102
rect 1840 2062 1880 2102
rect 1880 2062 1920 2102
rect 1920 2062 1960 2102
rect 1960 2062 2000 2102
rect 2000 2062 2040 2102
rect 2040 2062 2080 2102
rect 2080 2062 2120 2102
rect 2120 2062 2160 2102
rect 2160 2062 2200 2102
rect 2200 2062 2240 2102
rect 2240 2062 2280 2102
rect 2280 2062 2320 2102
rect 2320 2062 2360 2102
rect 2360 2062 2400 2102
rect 2400 2062 2440 2102
rect 2440 2062 2480 2102
rect 2480 2062 2520 2102
rect 2520 2062 2560 2102
rect 2560 2062 2600 2102
rect 2600 2062 2640 2102
rect 2640 2062 2680 2102
rect 2680 2062 2720 2102
rect 2720 2062 2760 2102
rect 2760 2062 2800 2102
rect 2800 2062 2840 2102
rect 2840 2062 2880 2102
rect 2880 2062 2920 2102
rect 2920 2062 2960 2102
rect 2960 2062 3000 2102
rect 3000 2062 3040 2102
rect 3040 2062 3080 2102
rect 3080 2062 3120 2102
rect 3120 2062 3160 2102
rect 3160 2062 3200 2102
rect 3200 2062 3240 2102
rect 3240 2062 3280 2102
rect 3280 2062 3320 2102
rect 3320 2062 3360 2102
rect 3360 2062 3400 2102
rect 3400 2062 3440 2102
rect 3440 2062 3480 2102
rect 3480 2062 3520 2102
rect 3520 2062 3560 2102
rect 3560 2062 3600 2102
rect 3600 2062 3640 2102
rect 3640 2062 3680 2102
rect 3680 2062 3720 2102
rect 3720 2062 3760 2102
rect 3760 2062 3800 2102
rect 3800 2062 3840 2102
rect 3840 2062 3880 2102
rect 3880 2062 3920 2102
rect 3920 2062 3960 2102
rect 3960 2062 4000 2102
rect 4000 2062 4040 2102
rect 4040 2062 4080 2102
rect 4080 2062 4120 2102
rect 4120 2062 4160 2102
rect 4160 2062 4200 2102
rect 4200 2062 4240 2102
rect 4240 2062 4280 2102
rect 16 79 56 119
rect 16 119 56 159
rect 16 159 56 199
rect 16 199 56 239
rect 16 239 56 279
rect 16 279 56 319
rect 16 319 56 359
rect 16 359 56 399
rect 16 399 56 439
rect 16 439 56 479
rect 16 479 56 519
rect 16 519 56 559
rect 16 559 56 599
rect 16 599 56 639
rect 16 639 56 679
rect 16 679 56 719
rect 16 719 56 759
rect 16 759 56 799
rect 16 799 56 839
rect 16 839 56 879
rect 16 879 56 919
rect 16 919 56 959
rect 16 959 56 999
rect 16 999 56 1039
rect 16 1039 56 1079
rect 16 1079 56 1119
rect 16 1119 56 1159
rect 16 1159 56 1199
rect 16 1199 56 1239
rect 16 1239 56 1279
rect 16 1279 56 1319
rect 16 1319 56 1359
rect 16 1359 56 1399
rect 16 1399 56 1439
rect 16 1439 56 1479
rect 16 1479 56 1519
rect 16 1519 56 1559
rect 16 1559 56 1599
rect 16 1599 56 1639
rect 16 1639 56 1679
rect 16 1679 56 1719
rect 16 1719 56 1759
rect 16 1759 56 1799
rect 16 1799 56 1839
rect 16 1839 56 1879
rect 16 1879 56 1919
rect 16 1919 56 1959
rect 16 1959 56 1999
rect 16 1999 56 2039
rect 4304 79 4344 119
rect 4304 119 4344 159
rect 4304 159 4344 199
rect 4304 199 4344 239
rect 4304 239 4344 279
rect 4304 279 4344 319
rect 4304 319 4344 359
rect 4304 359 4344 399
rect 4304 399 4344 439
rect 4304 439 4344 479
rect 4304 479 4344 519
rect 4304 519 4344 559
rect 4304 559 4344 599
rect 4304 599 4344 639
rect 4304 639 4344 679
rect 4304 679 4344 719
rect 4304 719 4344 759
rect 4304 759 4344 799
rect 4304 799 4344 839
rect 4304 839 4344 879
rect 4304 879 4344 919
rect 4304 919 4344 959
rect 4304 959 4344 999
rect 4304 999 4344 1039
rect 4304 1039 4344 1079
rect 4304 1079 4344 1119
rect 4304 1119 4344 1159
rect 4304 1159 4344 1199
rect 4304 1199 4344 1239
rect 4304 1239 4344 1279
rect 4304 1279 4344 1319
rect 4304 1319 4344 1359
rect 4304 1359 4344 1399
rect 4304 1399 4344 1439
rect 4304 1439 4344 1479
rect 4304 1479 4344 1519
rect 4304 1519 4344 1559
rect 4304 1559 4344 1599
rect 4304 1599 4344 1639
rect 4304 1639 4344 1679
rect 4304 1679 4344 1719
rect 4304 1719 4344 1759
rect 4304 1759 4344 1799
rect 4304 1799 4344 1839
rect 4304 1839 4344 1879
rect 4304 1879 4344 1919
rect 4304 1919 4344 1959
rect 4304 1959 4344 1999
rect 4304 1999 4344 2039
<< ptap >>
rect 0 0 4360 72
rect 0 2046 4360 2118
rect 0 0 72 2118
rect 4288 0 4360 2118
use JNWTR_RES16 XA1 
transform 1 0 344 0 1 344
box 344 344 4016 1774
<< labels >>
flabel locali s 8 8 4352 64 0 FreeSans 400 0 0 0 B
port 3 nsew signal bidirectional
flabel locali s 3764 1719 4052 1829 0 FreeSans 400 0 0 0 P
port 1 nsew signal bidirectional
flabel locali s 308 1719 596 1829 0 FreeSans 400 0 0 0 N
port 2 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 4360 2118
<< end >>
