

.subckt TGX2_CV A C B AVDD AVSS
MN0 AVSS C CN AVSS NCHDL
MN1 B C A AVSS NCHDL
MN1b B C A AVSS NCHDL

MP0 AVDD C CN AVDD PCHDL
MP1 B CN A AVDD PCHDL
MP1b B CN A AVDD PCHDL

.ends

.subckt DFTRIX1_CV D CK C CN Y AVDD AVSS
XA3 AVDD AVSS TAPCELLB_CV
XA2 D CK C NC QN AVDD AVSS DFRNQNX1_CV
XA0 QN C CN Y AVDD AVSS IVTRIX1_CV
.ends


.SUBCKT CKDIV2 AVDD AVSS CKI CKO CKO50DC RN
XA12v AVDD AVSS TAPCELLB_CV
XA1 CKI CKIB AVDD AVSS BFX1_CV
XA2 CKIB CKIN AVDD AVSS  IVX1_CV
XA4  QNI CKIN RN CKO50DC QN AVDD AVSS DFRNQNX1_CV
XA3 CKO50DC QNI AVDD AVSS  IVX1_CV
XA5 CKO50DC CKI CKO AVDD AVSS ANX1_CV
.ENDS

.subckt TOP AVDD AVSS
XA0 AVDD AVSS TAPCELLB_CV
XA1 Y1 AVDD AVSS TIEH_CV
XA2 Y2 AVDD AVSS TIEL_CV
XB0 AVDD AVSS TAPCELLB_CV
XB3 A3 Y3 AVDD AVSS IVX1_CV
XB4 A4 Y4 AVDD AVSS IVX2_CV
XB5 A5 Y5 AVDD AVSS IVX4_CV
XB6 A6 Y6 AVDD AVSS IVX8_CV
XC0 AVDD AVSS TAPCELLB_CV
XC7 A7 Y7 AVDD AVSS BFX1_CV
XD0 AVDD AVSS TAPCELLB_CV
XD8 A8 B8 Y8 AVDD AVSS NRX1_CV
XD9 A9 B9 Y9 AVDD AVSS NDX1_CV
XD10 A10 B10 Y10 AVDD AVSS ORX1_CV
XD11 A11 B11 Y11 AVDD AVSS ANX1_CV
XE0 AVDD AVSS TAPCELLB_CV
XE12 A12 Y12 AVDD AVSS SCX1_CV
XF0 AVDD AVSS TAPCELLB_CV
XF13 A13 Y13 V13 AVDD AVSS SWX2_CV
XF14 A14 Y14 V14 AVDD AVSS SWX4_CV
XF15 A15 Y15 V15 AVDD AVSS TGPD_CV
XG0 AVDD AVSS TAPCELLB_CV
XG1 A16 C16 B16 AVDD AVSS TGX2_CV
XH1 P17 N17 AVSS RPPO2 xoffset=4
XI1 P18 N18 AVSS RPPO4 xoffset=4
XJ1 P19 N19 AVSS RPPO8 xoffset=4
XK1 P20 N20 AVSS RPPO16 xoffset=4
XL0 AVDD AVSS TAPCELLB_CV xoffset=10
XL1 AVDD AVSS CKI21 CKO21 CKO50DC21 RN21 CKDIV2
XM0 AVDD AVSS TAPCELLB_CV
XM1 D22 CK22 C22 CN22 Y22 AVDD AVSS DFTRIX1_CV
XM2  D23 CK23 Q23 AVDD AVSS DFTSPCX1_CV
XN0 AVDD AVSS TAPCELLB_CV
XN1 A24 Y24  AVDD AVSS SCX1_CV
.ends
